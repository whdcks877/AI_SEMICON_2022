// Systolic Array
// JY Lee
// Version 2022-12-28

module SA
(
    input   wire                clk,
    input   wire                rst_n,

    //DATA part interface
    input   wire    [31:0]      data_i[24:0],   //temporary 32bit data, TODO: change size
    output  wire                dready_o,
    input   wire                dvalid_i,

    //Weight part interface
    input   wire    [31:0]      weight_i[399:0],    //temporary 32bit, 25X16 SA Matrix size
    input   wire                wvalid_i,
    output  wire                wready_o

    //accumulator interface
);
    reg     [31:0]      zero = 'd0;
    wire    [31:0]      data_o[24:0][15:0];
    wire    [31:0]      sum_o[24:0][15:0];

    //'0'th row
    PE u_pe0_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[0]),
        //Up part
        .weight_i(weight_i[0]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][0]),
        //Down part
        .sum_o(sum_o[0][0])
    );

    PE u_pe0_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][0]),
        //Up part
        .weight_i(weight_i[1]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][1]),
        //Down part
        .sum_o(sum_o[0][1])
    );

    PE u_pe0_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][1]),
        //Up part
        .weight_i(weight_i[2]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][2]),
        //Down part
        .sum_o(sum_o[0][2])
    );

    PE u_pe0_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][2]),
        //Up part
        .weight_i(weight_i[3]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][3]),
        //Down part
        .sum_o(sum_o[0][3])
    );

    PE u_pe0_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][3]),
        //Up part
        .weight_i(weight_i[4]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][4]),
        //Down part
        .sum_o(sum_o[0][4])
    );

    PE u_pe0_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][4]),
        //Up part
        .weight_i(weight_i[5]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][5]),
        //Down part
        .sum_o(sum_o[0][5])
    );

    PE u_pe0_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][5]),
        //Up part
        .weight_i(weight_i[6]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][6]),
        //Down part
        .sum_o(sum_o[0][6])
    );

    PE u_pe0_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][6]),
        //Up part
        .weight_i(weight_i[7]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][7]),
        //Down part
        .sum_o(sum_o[0][7])
    );

    PE u_pe0_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][7]),
        //Up part
        .weight_i(weight_i[8]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][8]),
        //Down part
        .sum_o(sum_o[0][8])
    );

    PE u_pe0_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][8]),
        //Up part
        .weight_i(weight_i[9]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][9]),
        //Down part
        .sum_o(sum_o[0][9])
    );

    PE u_pe0_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][9]),
        //Up part
        .weight_i(weight_i[10]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][10]),
        //Down part
        .sum_o(sum_o[0][10])
    );

    PE u_pe0_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][10]),
        //Up part
        .weight_i(weight_i[11]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][11]),
        //Down part
        .sum_o(sum_o[0][11])
    );

    PE u_pe0_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][11]),
        //Up part
        .weight_i(weight_i[12]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][12]),
        //Down part
        .sum_o(sum_o[0][12])
    );

    PE u_pe0_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][12]),
        //Up part
        .weight_i(weight_i[13]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][13]),
        //Down part
        .sum_o(sum_o[0][13])
    );

    PE u_pe0_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][13]),
        //Up part
        .weight_i(weight_i[14]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][14]),
        //Down part
        .sum_o(sum_o[0][14])
    );

    PE u_pe0_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[0][14]),
        //Up part
        .weight_i(weight_i[15]),
        .sum_i(zero),
        //Right part
        .data_o(data_o[0][15]),
        //Down part
        .sum_o(sum_o[0][15])
    );

    //'1'th row
    PE u_pe1_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[1]),
        //Up part
        .weight_i(weight_i[16]),
        .sum_i(sum_o[0][0]),
        //Right part
        .data_o(data_o[1][0]),
        //Down part
        .sum_o(sum_o[1][0])
    );

    PE u_pe1_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][0]),
        //Up part
        .weight_i(weight_i[17]),
        .sum_i(sum_o[0][1]),
        //Right part
        .data_o(data_o[1][1]),
        //Down part
        .sum_o(sum_o[1][1])
    );

    PE u_pe1_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][1]),
        //Up part
        .weight_i(weight_i[18]),
        .sum_i(sum_o[0][2]),
        //Right part
        .data_o(data_o[1][2]),
        //Down part
        .sum_o(sum_o[1][2])
    );

    PE u_pe1_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][2]),
        //Up part
        .weight_i(weight_i[19]),
        .sum_i(sum_o[0][3]),
        //Right part
        .data_o(data_o[1][3]),
        //Down part
        .sum_o(sum_o[1][3])
    );

    PE u_pe1_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][3]),
        //Up part
        .weight_i(weight_i[20]),
        .sum_i(sum_o[0][4]),
        //Right part
        .data_o(data_o[1][4]),
        //Down part
        .sum_o(sum_o[1][4])
    );

    PE u_pe1_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][4]),
        //Up part
        .weight_i(weight_i[21]),
        .sum_i(sum_o[0][5]),
        //Right part
        .data_o(data_o[1][5]),
        //Down part
        .sum_o(sum_o[1][5])
    );

    PE u_pe1_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][5]),
        //Up part
        .weight_i(weight_i[22]),
        .sum_i(sum_o[0][6]),
        //Right part
        .data_o(data_o[1][6]),
        //Down part
        .sum_o(sum_o[1][6])
    );

    PE u_pe1_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][6]),
        //Up part
        .weight_i(weight_i[23]),
        .sum_i(sum_o[0][7]),
        //Right part
        .data_o(data_o[1][7]),
        //Down part
        .sum_o(sum_o[1][7])
    );

    PE u_pe1_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][7]),
        //Up part
        .weight_i(weight_i[24]),
        .sum_i(sum_o[0][8]),
        //Right part
        .data_o(data_o[1][8]),
        //Down part
        .sum_o(sum_o[1][8])
    );

    PE u_pe1_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][8]),
        //Up part
        .weight_i(weight_i[25]),
        .sum_i(sum_o[0][9]),
        //Right part
        .data_o(data_o[1][9]),
        //Down part
        .sum_o(sum_o[1][9])
    );

    PE u_pe1_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][9]),
        //Up part
        .weight_i(weight_i[26]),
        .sum_i(sum_o[0][10]),
        //Right part
        .data_o(data_o[1][10]),
        //Down part
        .sum_o(sum_o[1][10])
    );

    PE u_pe1_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][10]),
        //Up part
        .weight_i(weight_i[27]),
        .sum_i(sum_o[0][11]),
        //Right part
        .data_o(data_o[1][11]),
        //Down part
        .sum_o(sum_o[1][11])
    );

    PE u_pe1_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][11]),
        //Up part
        .weight_i(weight_i[28]),
        .sum_i(sum_o[0][12]),
        //Right part
        .data_o(data_o[1][12]),
        //Down part
        .sum_o(sum_o[1][12])
    );

    PE u_pe1_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][12]),
        //Up part
        .weight_i(weight_i[29]),
        .sum_i(sum_o[0][13]),
        //Right part
        .data_o(data_o[1][13]),
        //Down part
        .sum_o(sum_o[1][13])
    );

    PE u_pe1_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][13]),
        //Up part
        .weight_i(weight_i[30]),
        .sum_i(sum_o[0][14]),
        //Right part
        .data_o(data_o[1][14]),
        //Down part
        .sum_o(sum_o[1][14])
    );

    PE u_pe1_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[1][14]),
        //Up part
        .weight_i(weight_i[31]),
        .sum_i(sum_o[0][15]),
        //Right part
        .data_o(data_o[1][15]),
        //Down part
        .sum_o(sum_o[1][15])
    );

    //'2'th row
    PE u_pe2_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[2]),
        //Up part
        .weight_i(weight_i[32]),
        .sum_i(sum_o[1][0]),
        //Right part
        .data_o(data_o[2][0]),
        //Down part
        .sum_o(sum_o[2][0])
    );

    PE u_pe2_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][0]),
        //Up part
        .weight_i(weight_i[33]),
        .sum_i(sum_o[1][1]),
        //Right part
        .data_o(data_o[2][1]),
        //Down part
        .sum_o(sum_o[2][1])
    );

    PE u_pe2_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][1]),
        //Up part
        .weight_i(weight_i[34]),
        .sum_i(sum_o[1][2]),
        //Right part
        .data_o(data_o[2][2]),
        //Down part
        .sum_o(sum_o[2][2])
    );

    PE u_pe2_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][2]),
        //Up part
        .weight_i(weight_i[35]),
        .sum_i(sum_o[1][3]),
        //Right part
        .data_o(data_o[2][3]),
        //Down part
        .sum_o(sum_o[2][3])
    );

    PE u_pe2_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][3]),
        //Up part
        .weight_i(weight_i[36]),
        .sum_i(sum_o[1][4]),
        //Right part
        .data_o(data_o[2][4]),
        //Down part
        .sum_o(sum_o[2][4])
    );

    PE u_pe2_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][4]),
        //Up part
        .weight_i(weight_i[37]),
        .sum_i(sum_o[1][5]),
        //Right part
        .data_o(data_o[2][5]),
        //Down part
        .sum_o(sum_o[2][5])
    );

    PE u_pe2_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][5]),
        //Up part
        .weight_i(weight_i[38]),
        .sum_i(sum_o[1][6]),
        //Right part
        .data_o(data_o[2][6]),
        //Down part
        .sum_o(sum_o[2][6])
    );

    PE u_pe2_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][6]),
        //Up part
        .weight_i(weight_i[39]),
        .sum_i(sum_o[1][7]),
        //Right part
        .data_o(data_o[2][7]),
        //Down part
        .sum_o(sum_o[2][7])
    );

    PE u_pe2_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][7]),
        //Up part
        .weight_i(weight_i[40]),
        .sum_i(sum_o[1][8]),
        //Right part
        .data_o(data_o[2][8]),
        //Down part
        .sum_o(sum_o[2][8])
    );

    PE u_pe2_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][8]),
        //Up part
        .weight_i(weight_i[41]),
        .sum_i(sum_o[1][9]),
        //Right part
        .data_o(data_o[2][9]),
        //Down part
        .sum_o(sum_o[2][9])
    );

    PE u_pe2_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][9]),
        //Up part
        .weight_i(weight_i[42]),
        .sum_i(sum_o[1][10]),
        //Right part
        .data_o(data_o[2][10]),
        //Down part
        .sum_o(sum_o[2][10])
    );

    PE u_pe2_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][10]),
        //Up part
        .weight_i(weight_i[43]),
        .sum_i(sum_o[1][11]),
        //Right part
        .data_o(data_o[2][11]),
        //Down part
        .sum_o(sum_o[2][11])
    );

    PE u_pe2_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][11]),
        //Up part
        .weight_i(weight_i[44]),
        .sum_i(sum_o[1][12]),
        //Right part
        .data_o(data_o[2][12]),
        //Down part
        .sum_o(sum_o[2][12])
    );

    PE u_pe2_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][12]),
        //Up part
        .weight_i(weight_i[45]),
        .sum_i(sum_o[1][13]),
        //Right part
        .data_o(data_o[2][13]),
        //Down part
        .sum_o(sum_o[2][13])
    );

    PE u_pe2_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][13]),
        //Up part
        .weight_i(weight_i[46]),
        .sum_i(sum_o[1][14]),
        //Right part
        .data_o(data_o[2][14]),
        //Down part
        .sum_o(sum_o[2][14])
    );

    PE u_pe2_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[2][14]),
        //Up part
        .weight_i(weight_i[47]),
        .sum_i(sum_o[1][15]),
        //Right part
        .data_o(data_o[2][15]),
        //Down part
        .sum_o(sum_o[2][15])
    );

    //'3'th row
    PE u_pe3_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[3]),
        //Up part
        .weight_i(weight_i[48]),
        .sum_i(sum_o[2][0]),
        //Right part
        .data_o(data_o[3][0]),
        //Down part
        .sum_o(sum_o[3][0])
    );

    PE u_pe3_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][0]),
        //Up part
        .weight_i(weight_i[49]),
        .sum_i(sum_o[2][1]),
        //Right part
        .data_o(data_o[3][1]),
        //Down part
        .sum_o(sum_o[3][1])
    );

    PE u_pe3_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][1]),
        //Up part
        .weight_i(weight_i[50]),
        .sum_i(sum_o[2][2]),
        //Right part
        .data_o(data_o[3][2]),
        //Down part
        .sum_o(sum_o[3][2])
    );

    PE u_pe3_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][2]),
        //Up part
        .weight_i(weight_i[51]),
        .sum_i(sum_o[2][3]),
        //Right part
        .data_o(data_o[3][3]),
        //Down part
        .sum_o(sum_o[3][3])
    );

    PE u_pe3_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][3]),
        //Up part
        .weight_i(weight_i[52]),
        .sum_i(sum_o[2][4]),
        //Right part
        .data_o(data_o[3][4]),
        //Down part
        .sum_o(sum_o[3][4])
    );

    PE u_pe3_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][4]),
        //Up part
        .weight_i(weight_i[53]),
        .sum_i(sum_o[2][5]),
        //Right part
        .data_o(data_o[3][5]),
        //Down part
        .sum_o(sum_o[3][5])
    );

    PE u_pe3_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][5]),
        //Up part
        .weight_i(weight_i[54]),
        .sum_i(sum_o[2][6]),
        //Right part
        .data_o(data_o[3][6]),
        //Down part
        .sum_o(sum_o[3][6])
    );

    PE u_pe3_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][6]),
        //Up part
        .weight_i(weight_i[55]),
        .sum_i(sum_o[2][7]),
        //Right part
        .data_o(data_o[3][7]),
        //Down part
        .sum_o(sum_o[3][7])
    );

    PE u_pe3_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][7]),
        //Up part
        .weight_i(weight_i[56]),
        .sum_i(sum_o[2][8]),
        //Right part
        .data_o(data_o[3][8]),
        //Down part
        .sum_o(sum_o[3][8])
    );

    PE u_pe3_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][8]),
        //Up part
        .weight_i(weight_i[57]),
        .sum_i(sum_o[2][9]),
        //Right part
        .data_o(data_o[3][9]),
        //Down part
        .sum_o(sum_o[3][9])
    );

    PE u_pe3_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][9]),
        //Up part
        .weight_i(weight_i[58]),
        .sum_i(sum_o[2][10]),
        //Right part
        .data_o(data_o[3][10]),
        //Down part
        .sum_o(sum_o[3][10])
    );

    PE u_pe3_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][10]),
        //Up part
        .weight_i(weight_i[59]),
        .sum_i(sum_o[2][11]),
        //Right part
        .data_o(data_o[3][11]),
        //Down part
        .sum_o(sum_o[3][11])
    );

    PE u_pe3_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][11]),
        //Up part
        .weight_i(weight_i[60]),
        .sum_i(sum_o[2][12]),
        //Right part
        .data_o(data_o[3][12]),
        //Down part
        .sum_o(sum_o[3][12])
    );

    PE u_pe3_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][12]),
        //Up part
        .weight_i(weight_i[61]),
        .sum_i(sum_o[2][13]),
        //Right part
        .data_o(data_o[3][13]),
        //Down part
        .sum_o(sum_o[3][13])
    );

    PE u_pe3_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][13]),
        //Up part
        .weight_i(weight_i[62]),
        .sum_i(sum_o[2][14]),
        //Right part
        .data_o(data_o[3][14]),
        //Down part
        .sum_o(sum_o[3][14])
    );

    PE u_pe3_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[3][14]),
        //Up part
        .weight_i(weight_i[63]),
        .sum_i(sum_o[2][15]),
        //Right part
        .data_o(data_o[3][15]),
        //Down part
        .sum_o(sum_o[3][15])
    );

    //'4'th row
    PE u_pe4_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[4]),
        //Up part
        .weight_i(weight_i[64]),
        .sum_i(sum_o[3][0]),
        //Right part
        .data_o(data_o[4][0]),
        //Down part
        .sum_o(sum_o[4][0])
    );

    PE u_pe4_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][0]),
        //Up part
        .weight_i(weight_i[65]),
        .sum_i(sum_o[3][1]),
        //Right part
        .data_o(data_o[4][1]),
        //Down part
        .sum_o(sum_o[4][1])
    );

    PE u_pe4_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][1]),
        //Up part
        .weight_i(weight_i[66]),
        .sum_i(sum_o[3][2]),
        //Right part
        .data_o(data_o[4][2]),
        //Down part
        .sum_o(sum_o[4][2])
    );

    PE u_pe4_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][2]),
        //Up part
        .weight_i(weight_i[67]),
        .sum_i(sum_o[3][3]),
        //Right part
        .data_o(data_o[4][3]),
        //Down part
        .sum_o(sum_o[4][3])
    );

    PE u_pe4_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][3]),
        //Up part
        .weight_i(weight_i[68]),
        .sum_i(sum_o[3][4]),
        //Right part
        .data_o(data_o[4][4]),
        //Down part
        .sum_o(sum_o[4][4])
    );

    PE u_pe4_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][4]),
        //Up part
        .weight_i(weight_i[69]),
        .sum_i(sum_o[3][5]),
        //Right part
        .data_o(data_o[4][5]),
        //Down part
        .sum_o(sum_o[4][5])
    );

    PE u_pe4_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][5]),
        //Up part
        .weight_i(weight_i[70]),
        .sum_i(sum_o[3][6]),
        //Right part
        .data_o(data_o[4][6]),
        //Down part
        .sum_o(sum_o[4][6])
    );

    PE u_pe4_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][6]),
        //Up part
        .weight_i(weight_i[71]),
        .sum_i(sum_o[3][7]),
        //Right part
        .data_o(data_o[4][7]),
        //Down part
        .sum_o(sum_o[4][7])
    );

    PE u_pe4_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][7]),
        //Up part
        .weight_i(weight_i[72]),
        .sum_i(sum_o[3][8]),
        //Right part
        .data_o(data_o[4][8]),
        //Down part
        .sum_o(sum_o[4][8])
    );

    PE u_pe4_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][8]),
        //Up part
        .weight_i(weight_i[73]),
        .sum_i(sum_o[3][9]),
        //Right part
        .data_o(data_o[4][9]),
        //Down part
        .sum_o(sum_o[4][9])
    );

    PE u_pe4_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][9]),
        //Up part
        .weight_i(weight_i[74]),
        .sum_i(sum_o[3][10]),
        //Right part
        .data_o(data_o[4][10]),
        //Down part
        .sum_o(sum_o[4][10])
    );

    PE u_pe4_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][10]),
        //Up part
        .weight_i(weight_i[75]),
        .sum_i(sum_o[3][11]),
        //Right part
        .data_o(data_o[4][11]),
        //Down part
        .sum_o(sum_o[4][11])
    );

    PE u_pe4_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][11]),
        //Up part
        .weight_i(weight_i[76]),
        .sum_i(sum_o[3][12]),
        //Right part
        .data_o(data_o[4][12]),
        //Down part
        .sum_o(sum_o[4][12])
    );

    PE u_pe4_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][12]),
        //Up part
        .weight_i(weight_i[77]),
        .sum_i(sum_o[3][13]),
        //Right part
        .data_o(data_o[4][13]),
        //Down part
        .sum_o(sum_o[4][13])
    );

    PE u_pe4_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][13]),
        //Up part
        .weight_i(weight_i[78]),
        .sum_i(sum_o[3][14]),
        //Right part
        .data_o(data_o[4][14]),
        //Down part
        .sum_o(sum_o[4][14])
    );

    PE u_pe4_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[4][14]),
        //Up part
        .weight_i(weight_i[79]),
        .sum_i(sum_o[3][15]),
        //Right part
        .data_o(data_o[4][15]),
        //Down part
        .sum_o(sum_o[4][15])
    );

    //'5'th row
    PE u_pe5_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[5]),
        //Up part
        .weight_i(weight_i[80]),
        .sum_i(sum_o[4][0]),
        //Right part
        .data_o(data_o[5][0]),
        //Down part
        .sum_o(sum_o[5][0])
    );

    PE u_pe5_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][0]),
        //Up part
        .weight_i(weight_i[81]),
        .sum_i(sum_o[4][1]),
        //Right part
        .data_o(data_o[5][1]),
        //Down part
        .sum_o(sum_o[5][1])
    );

    PE u_pe5_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][1]),
        //Up part
        .weight_i(weight_i[82]),
        .sum_i(sum_o[4][2]),
        //Right part
        .data_o(data_o[5][2]),
        //Down part
        .sum_o(sum_o[5][2])
    );

    PE u_pe5_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][2]),
        //Up part
        .weight_i(weight_i[83]),
        .sum_i(sum_o[4][3]),
        //Right part
        .data_o(data_o[5][3]),
        //Down part
        .sum_o(sum_o[5][3])
    );

    PE u_pe5_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][3]),
        //Up part
        .weight_i(weight_i[84]),
        .sum_i(sum_o[4][4]),
        //Right part
        .data_o(data_o[5][4]),
        //Down part
        .sum_o(sum_o[5][4])
    );

    PE u_pe5_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][4]),
        //Up part
        .weight_i(weight_i[85]),
        .sum_i(sum_o[4][5]),
        //Right part
        .data_o(data_o[5][5]),
        //Down part
        .sum_o(sum_o[5][5])
    );

    PE u_pe5_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][5]),
        //Up part
        .weight_i(weight_i[86]),
        .sum_i(sum_o[4][6]),
        //Right part
        .data_o(data_o[5][6]),
        //Down part
        .sum_o(sum_o[5][6])
    );

    PE u_pe5_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][6]),
        //Up part
        .weight_i(weight_i[87]),
        .sum_i(sum_o[4][7]),
        //Right part
        .data_o(data_o[5][7]),
        //Down part
        .sum_o(sum_o[5][7])
    );

    PE u_pe5_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][7]),
        //Up part
        .weight_i(weight_i[88]),
        .sum_i(sum_o[4][8]),
        //Right part
        .data_o(data_o[5][8]),
        //Down part
        .sum_o(sum_o[5][8])
    );

    PE u_pe5_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][8]),
        //Up part
        .weight_i(weight_i[89]),
        .sum_i(sum_o[4][9]),
        //Right part
        .data_o(data_o[5][9]),
        //Down part
        .sum_o(sum_o[5][9])
    );

    PE u_pe5_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][9]),
        //Up part
        .weight_i(weight_i[90]),
        .sum_i(sum_o[4][10]),
        //Right part
        .data_o(data_o[5][10]),
        //Down part
        .sum_o(sum_o[5][10])
    );

    PE u_pe5_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][10]),
        //Up part
        .weight_i(weight_i[91]),
        .sum_i(sum_o[4][11]),
        //Right part
        .data_o(data_o[5][11]),
        //Down part
        .sum_o(sum_o[5][11])
    );

    PE u_pe5_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][11]),
        //Up part
        .weight_i(weight_i[92]),
        .sum_i(sum_o[4][12]),
        //Right part
        .data_o(data_o[5][12]),
        //Down part
        .sum_o(sum_o[5][12])
    );

    PE u_pe5_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][12]),
        //Up part
        .weight_i(weight_i[93]),
        .sum_i(sum_o[4][13]),
        //Right part
        .data_o(data_o[5][13]),
        //Down part
        .sum_o(sum_o[5][13])
    );

    PE u_pe5_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][13]),
        //Up part
        .weight_i(weight_i[94]),
        .sum_i(sum_o[4][14]),
        //Right part
        .data_o(data_o[5][14]),
        //Down part
        .sum_o(sum_o[5][14])
    );

    PE u_pe5_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[5][14]),
        //Up part
        .weight_i(weight_i[95]),
        .sum_i(sum_o[4][15]),
        //Right part
        .data_o(data_o[5][15]),
        //Down part
        .sum_o(sum_o[5][15])
    );

    //'6'th row
    PE u_pe6_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[6]),
        //Up part
        .weight_i(weight_i[96]),
        .sum_i(sum_o[5][0]),
        //Right part
        .data_o(data_o[6][0]),
        //Down part
        .sum_o(sum_o[6][0])
    );

    PE u_pe6_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][0]),
        //Up part
        .weight_i(weight_i[97]),
        .sum_i(sum_o[5][1]),
        //Right part
        .data_o(data_o[6][1]),
        //Down part
        .sum_o(sum_o[6][1])
    );

    PE u_pe6_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][1]),
        //Up part
        .weight_i(weight_i[98]),
        .sum_i(sum_o[5][2]),
        //Right part
        .data_o(data_o[6][2]),
        //Down part
        .sum_o(sum_o[6][2])
    );

    PE u_pe6_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][2]),
        //Up part
        .weight_i(weight_i[99]),
        .sum_i(sum_o[5][3]),
        //Right part
        .data_o(data_o[6][3]),
        //Down part
        .sum_o(sum_o[6][3])
    );

    PE u_pe6_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][3]),
        //Up part
        .weight_i(weight_i[100]),
        .sum_i(sum_o[5][4]),
        //Right part
        .data_o(data_o[6][4]),
        //Down part
        .sum_o(sum_o[6][4])
    );

    PE u_pe6_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][4]),
        //Up part
        .weight_i(weight_i[101]),
        .sum_i(sum_o[5][5]),
        //Right part
        .data_o(data_o[6][5]),
        //Down part
        .sum_o(sum_o[6][5])
    );

    PE u_pe6_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][5]),
        //Up part
        .weight_i(weight_i[102]),
        .sum_i(sum_o[5][6]),
        //Right part
        .data_o(data_o[6][6]),
        //Down part
        .sum_o(sum_o[6][6])
    );

    PE u_pe6_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][6]),
        //Up part
        .weight_i(weight_i[103]),
        .sum_i(sum_o[5][7]),
        //Right part
        .data_o(data_o[6][7]),
        //Down part
        .sum_o(sum_o[6][7])
    );

    PE u_pe6_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][7]),
        //Up part
        .weight_i(weight_i[104]),
        .sum_i(sum_o[5][8]),
        //Right part
        .data_o(data_o[6][8]),
        //Down part
        .sum_o(sum_o[6][8])
    );

    PE u_pe6_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][8]),
        //Up part
        .weight_i(weight_i[105]),
        .sum_i(sum_o[5][9]),
        //Right part
        .data_o(data_o[6][9]),
        //Down part
        .sum_o(sum_o[6][9])
    );

    PE u_pe6_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][9]),
        //Up part
        .weight_i(weight_i[106]),
        .sum_i(sum_o[5][10]),
        //Right part
        .data_o(data_o[6][10]),
        //Down part
        .sum_o(sum_o[6][10])
    );

    PE u_pe6_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][10]),
        //Up part
        .weight_i(weight_i[107]),
        .sum_i(sum_o[5][11]),
        //Right part
        .data_o(data_o[6][11]),
        //Down part
        .sum_o(sum_o[6][11])
    );

    PE u_pe6_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][11]),
        //Up part
        .weight_i(weight_i[108]),
        .sum_i(sum_o[5][12]),
        //Right part
        .data_o(data_o[6][12]),
        //Down part
        .sum_o(sum_o[6][12])
    );

    PE u_pe6_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][12]),
        //Up part
        .weight_i(weight_i[109]),
        .sum_i(sum_o[5][13]),
        //Right part
        .data_o(data_o[6][13]),
        //Down part
        .sum_o(sum_o[6][13])
    );

    PE u_pe6_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][13]),
        //Up part
        .weight_i(weight_i[110]),
        .sum_i(sum_o[5][14]),
        //Right part
        .data_o(data_o[6][14]),
        //Down part
        .sum_o(sum_o[6][14])
    );

    PE u_pe6_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[6][14]),
        //Up part
        .weight_i(weight_i[111]),
        .sum_i(sum_o[5][15]),
        //Right part
        .data_o(data_o[6][15]),
        //Down part
        .sum_o(sum_o[6][15])
    );

    //'7'th row
    PE u_pe7_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[7]),
        //Up part
        .weight_i(weight_i[112]),
        .sum_i(sum_o[6][0]),
        //Right part
        .data_o(data_o[7][0]),
        //Down part
        .sum_o(sum_o[7][0])
    );

    PE u_pe7_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][0]),
        //Up part
        .weight_i(weight_i[113]),
        .sum_i(sum_o[6][1]),
        //Right part
        .data_o(data_o[7][1]),
        //Down part
        .sum_o(sum_o[7][1])
    );

    PE u_pe7_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][1]),
        //Up part
        .weight_i(weight_i[114]),
        .sum_i(sum_o[6][2]),
        //Right part
        .data_o(data_o[7][2]),
        //Down part
        .sum_o(sum_o[7][2])
    );

    PE u_pe7_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][2]),
        //Up part
        .weight_i(weight_i[115]),
        .sum_i(sum_o[6][3]),
        //Right part
        .data_o(data_o[7][3]),
        //Down part
        .sum_o(sum_o[7][3])
    );

    PE u_pe7_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][3]),
        //Up part
        .weight_i(weight_i[116]),
        .sum_i(sum_o[6][4]),
        //Right part
        .data_o(data_o[7][4]),
        //Down part
        .sum_o(sum_o[7][4])
    );

    PE u_pe7_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][4]),
        //Up part
        .weight_i(weight_i[117]),
        .sum_i(sum_o[6][5]),
        //Right part
        .data_o(data_o[7][5]),
        //Down part
        .sum_o(sum_o[7][5])
    );

    PE u_pe7_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][5]),
        //Up part
        .weight_i(weight_i[118]),
        .sum_i(sum_o[6][6]),
        //Right part
        .data_o(data_o[7][6]),
        //Down part
        .sum_o(sum_o[7][6])
    );

    PE u_pe7_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][6]),
        //Up part
        .weight_i(weight_i[119]),
        .sum_i(sum_o[6][7]),
        //Right part
        .data_o(data_o[7][7]),
        //Down part
        .sum_o(sum_o[7][7])
    );

    PE u_pe7_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][7]),
        //Up part
        .weight_i(weight_i[120]),
        .sum_i(sum_o[6][8]),
        //Right part
        .data_o(data_o[7][8]),
        //Down part
        .sum_o(sum_o[7][8])
    );

    PE u_pe7_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][8]),
        //Up part
        .weight_i(weight_i[121]),
        .sum_i(sum_o[6][9]),
        //Right part
        .data_o(data_o[7][9]),
        //Down part
        .sum_o(sum_o[7][9])
    );

    PE u_pe7_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][9]),
        //Up part
        .weight_i(weight_i[122]),
        .sum_i(sum_o[6][10]),
        //Right part
        .data_o(data_o[7][10]),
        //Down part
        .sum_o(sum_o[7][10])
    );

    PE u_pe7_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][10]),
        //Up part
        .weight_i(weight_i[123]),
        .sum_i(sum_o[6][11]),
        //Right part
        .data_o(data_o[7][11]),
        //Down part
        .sum_o(sum_o[7][11])
    );

    PE u_pe7_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][11]),
        //Up part
        .weight_i(weight_i[124]),
        .sum_i(sum_o[6][12]),
        //Right part
        .data_o(data_o[7][12]),
        //Down part
        .sum_o(sum_o[7][12])
    );

    PE u_pe7_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][12]),
        //Up part
        .weight_i(weight_i[125]),
        .sum_i(sum_o[6][13]),
        //Right part
        .data_o(data_o[7][13]),
        //Down part
        .sum_o(sum_o[7][13])
    );

    PE u_pe7_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][13]),
        //Up part
        .weight_i(weight_i[126]),
        .sum_i(sum_o[6][14]),
        //Right part
        .data_o(data_o[7][14]),
        //Down part
        .sum_o(sum_o[7][14])
    );

    PE u_pe7_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[7][14]),
        //Up part
        .weight_i(weight_i[127]),
        .sum_i(sum_o[6][15]),
        //Right part
        .data_o(data_o[7][15]),
        //Down part
        .sum_o(sum_o[7][15])
    );

    //'8'th row
    PE u_pe8_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[8]),
        //Up part
        .weight_i(weight_i[128]),
        .sum_i(sum_o[7][0]),
        //Right part
        .data_o(data_o[8][0]),
        //Down part
        .sum_o(sum_o[8][0])
    );

    PE u_pe8_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][0]),
        //Up part
        .weight_i(weight_i[129]),
        .sum_i(sum_o[7][1]),
        //Right part
        .data_o(data_o[8][1]),
        //Down part
        .sum_o(sum_o[8][1])
    );

    PE u_pe8_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][1]),
        //Up part
        .weight_i(weight_i[130]),
        .sum_i(sum_o[7][2]),
        //Right part
        .data_o(data_o[8][2]),
        //Down part
        .sum_o(sum_o[8][2])
    );

    PE u_pe8_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][2]),
        //Up part
        .weight_i(weight_i[131]),
        .sum_i(sum_o[7][3]),
        //Right part
        .data_o(data_o[8][3]),
        //Down part
        .sum_o(sum_o[8][3])
    );

    PE u_pe8_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][3]),
        //Up part
        .weight_i(weight_i[132]),
        .sum_i(sum_o[7][4]),
        //Right part
        .data_o(data_o[8][4]),
        //Down part
        .sum_o(sum_o[8][4])
    );

    PE u_pe8_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][4]),
        //Up part
        .weight_i(weight_i[133]),
        .sum_i(sum_o[7][5]),
        //Right part
        .data_o(data_o[8][5]),
        //Down part
        .sum_o(sum_o[8][5])
    );

    PE u_pe8_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][5]),
        //Up part
        .weight_i(weight_i[134]),
        .sum_i(sum_o[7][6]),
        //Right part
        .data_o(data_o[8][6]),
        //Down part
        .sum_o(sum_o[8][6])
    );

    PE u_pe8_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][6]),
        //Up part
        .weight_i(weight_i[135]),
        .sum_i(sum_o[7][7]),
        //Right part
        .data_o(data_o[8][7]),
        //Down part
        .sum_o(sum_o[8][7])
    );

    PE u_pe8_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][7]),
        //Up part
        .weight_i(weight_i[136]),
        .sum_i(sum_o[7][8]),
        //Right part
        .data_o(data_o[8][8]),
        //Down part
        .sum_o(sum_o[8][8])
    );

    PE u_pe8_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][8]),
        //Up part
        .weight_i(weight_i[137]),
        .sum_i(sum_o[7][9]),
        //Right part
        .data_o(data_o[8][9]),
        //Down part
        .sum_o(sum_o[8][9])
    );

    PE u_pe8_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][9]),
        //Up part
        .weight_i(weight_i[138]),
        .sum_i(sum_o[7][10]),
        //Right part
        .data_o(data_o[8][10]),
        //Down part
        .sum_o(sum_o[8][10])
    );

    PE u_pe8_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][10]),
        //Up part
        .weight_i(weight_i[139]),
        .sum_i(sum_o[7][11]),
        //Right part
        .data_o(data_o[8][11]),
        //Down part
        .sum_o(sum_o[8][11])
    );

    PE u_pe8_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][11]),
        //Up part
        .weight_i(weight_i[140]),
        .sum_i(sum_o[7][12]),
        //Right part
        .data_o(data_o[8][12]),
        //Down part
        .sum_o(sum_o[8][12])
    );

    PE u_pe8_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][12]),
        //Up part
        .weight_i(weight_i[141]),
        .sum_i(sum_o[7][13]),
        //Right part
        .data_o(data_o[8][13]),
        //Down part
        .sum_o(sum_o[8][13])
    );

    PE u_pe8_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][13]),
        //Up part
        .weight_i(weight_i[142]),
        .sum_i(sum_o[7][14]),
        //Right part
        .data_o(data_o[8][14]),
        //Down part
        .sum_o(sum_o[8][14])
    );

    PE u_pe8_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[8][14]),
        //Up part
        .weight_i(weight_i[143]),
        .sum_i(sum_o[7][15]),
        //Right part
        .data_o(data_o[8][15]),
        //Down part
        .sum_o(sum_o[8][15])
    );

    //'9'th row
    PE u_pe9_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[9]),
        //Up part
        .weight_i(weight_i[144]),
        .sum_i(sum_o[8][0]),
        //Right part
        .data_o(data_o[9][0]),
        //Down part
        .sum_o(sum_o[9][0])
    );

    PE u_pe9_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][0]),
        //Up part
        .weight_i(weight_i[145]),
        .sum_i(sum_o[8][1]),
        //Right part
        .data_o(data_o[9][1]),
        //Down part
        .sum_o(sum_o[9][1])
    );

    PE u_pe9_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][1]),
        //Up part
        .weight_i(weight_i[146]),
        .sum_i(sum_o[8][2]),
        //Right part
        .data_o(data_o[9][2]),
        //Down part
        .sum_o(sum_o[9][2])
    );

    PE u_pe9_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][2]),
        //Up part
        .weight_i(weight_i[147]),
        .sum_i(sum_o[8][3]),
        //Right part
        .data_o(data_o[9][3]),
        //Down part
        .sum_o(sum_o[9][3])
    );

    PE u_pe9_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][3]),
        //Up part
        .weight_i(weight_i[148]),
        .sum_i(sum_o[8][4]),
        //Right part
        .data_o(data_o[9][4]),
        //Down part
        .sum_o(sum_o[9][4])
    );

    PE u_pe9_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][4]),
        //Up part
        .weight_i(weight_i[149]),
        .sum_i(sum_o[8][5]),
        //Right part
        .data_o(data_o[9][5]),
        //Down part
        .sum_o(sum_o[9][5])
    );

    PE u_pe9_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][5]),
        //Up part
        .weight_i(weight_i[150]),
        .sum_i(sum_o[8][6]),
        //Right part
        .data_o(data_o[9][6]),
        //Down part
        .sum_o(sum_o[9][6])
    );

    PE u_pe9_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][6]),
        //Up part
        .weight_i(weight_i[151]),
        .sum_i(sum_o[8][7]),
        //Right part
        .data_o(data_o[9][7]),
        //Down part
        .sum_o(sum_o[9][7])
    );

    PE u_pe9_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][7]),
        //Up part
        .weight_i(weight_i[152]),
        .sum_i(sum_o[8][8]),
        //Right part
        .data_o(data_o[9][8]),
        //Down part
        .sum_o(sum_o[9][8])
    );

    PE u_pe9_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][8]),
        //Up part
        .weight_i(weight_i[153]),
        .sum_i(sum_o[8][9]),
        //Right part
        .data_o(data_o[9][9]),
        //Down part
        .sum_o(sum_o[9][9])
    );

    PE u_pe9_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][9]),
        //Up part
        .weight_i(weight_i[154]),
        .sum_i(sum_o[8][10]),
        //Right part
        .data_o(data_o[9][10]),
        //Down part
        .sum_o(sum_o[9][10])
    );

    PE u_pe9_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][10]),
        //Up part
        .weight_i(weight_i[155]),
        .sum_i(sum_o[8][11]),
        //Right part
        .data_o(data_o[9][11]),
        //Down part
        .sum_o(sum_o[9][11])
    );

    PE u_pe9_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][11]),
        //Up part
        .weight_i(weight_i[156]),
        .sum_i(sum_o[8][12]),
        //Right part
        .data_o(data_o[9][12]),
        //Down part
        .sum_o(sum_o[9][12])
    );

    PE u_pe9_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][12]),
        //Up part
        .weight_i(weight_i[157]),
        .sum_i(sum_o[8][13]),
        //Right part
        .data_o(data_o[9][13]),
        //Down part
        .sum_o(sum_o[9][13])
    );

    PE u_pe9_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][13]),
        //Up part
        .weight_i(weight_i[158]),
        .sum_i(sum_o[8][14]),
        //Right part
        .data_o(data_o[9][14]),
        //Down part
        .sum_o(sum_o[9][14])
    );

    PE u_pe9_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[9][14]),
        //Up part
        .weight_i(weight_i[159]),
        .sum_i(sum_o[8][15]),
        //Right part
        .data_o(data_o[9][15]),
        //Down part
        .sum_o(sum_o[9][15])
    );

    //'10'th row
    PE u_pe10_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[10]),
        //Up part
        .weight_i(weight_i[160]),
        .sum_i(sum_o[9][0]),
        //Right part
        .data_o(data_o[10][0]),
        //Down part
        .sum_o(sum_o[10][0])
    );

    PE u_pe10_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][0]),
        //Up part
        .weight_i(weight_i[161]),
        .sum_i(sum_o[9][1]),
        //Right part
        .data_o(data_o[10][1]),
        //Down part
        .sum_o(sum_o[10][1])
    );

    PE u_pe10_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][1]),
        //Up part
        .weight_i(weight_i[162]),
        .sum_i(sum_o[9][2]),
        //Right part
        .data_o(data_o[10][2]),
        //Down part
        .sum_o(sum_o[10][2])
    );

    PE u_pe10_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][2]),
        //Up part
        .weight_i(weight_i[163]),
        .sum_i(sum_o[9][3]),
        //Right part
        .data_o(data_o[10][3]),
        //Down part
        .sum_o(sum_o[10][3])
    );

    PE u_pe10_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][3]),
        //Up part
        .weight_i(weight_i[164]),
        .sum_i(sum_o[9][4]),
        //Right part
        .data_o(data_o[10][4]),
        //Down part
        .sum_o(sum_o[10][4])
    );

    PE u_pe10_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][4]),
        //Up part
        .weight_i(weight_i[165]),
        .sum_i(sum_o[9][5]),
        //Right part
        .data_o(data_o[10][5]),
        //Down part
        .sum_o(sum_o[10][5])
    );

    PE u_pe10_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][5]),
        //Up part
        .weight_i(weight_i[166]),
        .sum_i(sum_o[9][6]),
        //Right part
        .data_o(data_o[10][6]),
        //Down part
        .sum_o(sum_o[10][6])
    );

    PE u_pe10_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][6]),
        //Up part
        .weight_i(weight_i[167]),
        .sum_i(sum_o[9][7]),
        //Right part
        .data_o(data_o[10][7]),
        //Down part
        .sum_o(sum_o[10][7])
    );

    PE u_pe10_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][7]),
        //Up part
        .weight_i(weight_i[168]),
        .sum_i(sum_o[9][8]),
        //Right part
        .data_o(data_o[10][8]),
        //Down part
        .sum_o(sum_o[10][8])
    );

    PE u_pe10_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][8]),
        //Up part
        .weight_i(weight_i[169]),
        .sum_i(sum_o[9][9]),
        //Right part
        .data_o(data_o[10][9]),
        //Down part
        .sum_o(sum_o[10][9])
    );

    PE u_pe10_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][9]),
        //Up part
        .weight_i(weight_i[170]),
        .sum_i(sum_o[9][10]),
        //Right part
        .data_o(data_o[10][10]),
        //Down part
        .sum_o(sum_o[10][10])
    );

    PE u_pe10_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][10]),
        //Up part
        .weight_i(weight_i[171]),
        .sum_i(sum_o[9][11]),
        //Right part
        .data_o(data_o[10][11]),
        //Down part
        .sum_o(sum_o[10][11])
    );

    PE u_pe10_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][11]),
        //Up part
        .weight_i(weight_i[172]),
        .sum_i(sum_o[9][12]),
        //Right part
        .data_o(data_o[10][12]),
        //Down part
        .sum_o(sum_o[10][12])
    );

    PE u_pe10_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][12]),
        //Up part
        .weight_i(weight_i[173]),
        .sum_i(sum_o[9][13]),
        //Right part
        .data_o(data_o[10][13]),
        //Down part
        .sum_o(sum_o[10][13])
    );

    PE u_pe10_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][13]),
        //Up part
        .weight_i(weight_i[174]),
        .sum_i(sum_o[9][14]),
        //Right part
        .data_o(data_o[10][14]),
        //Down part
        .sum_o(sum_o[10][14])
    );

    PE u_pe10_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[10][14]),
        //Up part
        .weight_i(weight_i[175]),
        .sum_i(sum_o[9][15]),
        //Right part
        .data_o(data_o[10][15]),
        //Down part
        .sum_o(sum_o[10][15])
    );

    //'11'th row
    PE u_pe11_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[11]),
        //Up part
        .weight_i(weight_i[176]),
        .sum_i(sum_o[10][0]),
        //Right part
        .data_o(data_o[11][0]),
        //Down part
        .sum_o(sum_o[11][0])
    );

    PE u_pe11_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][0]),
        //Up part
        .weight_i(weight_i[177]),
        .sum_i(sum_o[10][1]),
        //Right part
        .data_o(data_o[11][1]),
        //Down part
        .sum_o(sum_o[11][1])
    );

    PE u_pe11_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][1]),
        //Up part
        .weight_i(weight_i[178]),
        .sum_i(sum_o[10][2]),
        //Right part
        .data_o(data_o[11][2]),
        //Down part
        .sum_o(sum_o[11][2])
    );

    PE u_pe11_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][2]),
        //Up part
        .weight_i(weight_i[179]),
        .sum_i(sum_o[10][3]),
        //Right part
        .data_o(data_o[11][3]),
        //Down part
        .sum_o(sum_o[11][3])
    );

    PE u_pe11_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][3]),
        //Up part
        .weight_i(weight_i[180]),
        .sum_i(sum_o[10][4]),
        //Right part
        .data_o(data_o[11][4]),
        //Down part
        .sum_o(sum_o[11][4])
    );

    PE u_pe11_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][4]),
        //Up part
        .weight_i(weight_i[181]),
        .sum_i(sum_o[10][5]),
        //Right part
        .data_o(data_o[11][5]),
        //Down part
        .sum_o(sum_o[11][5])
    );

    PE u_pe11_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][5]),
        //Up part
        .weight_i(weight_i[182]),
        .sum_i(sum_o[10][6]),
        //Right part
        .data_o(data_o[11][6]),
        //Down part
        .sum_o(sum_o[11][6])
    );

    PE u_pe11_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][6]),
        //Up part
        .weight_i(weight_i[183]),
        .sum_i(sum_o[10][7]),
        //Right part
        .data_o(data_o[11][7]),
        //Down part
        .sum_o(sum_o[11][7])
    );

    PE u_pe11_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][7]),
        //Up part
        .weight_i(weight_i[184]),
        .sum_i(sum_o[10][8]),
        //Right part
        .data_o(data_o[11][8]),
        //Down part
        .sum_o(sum_o[11][8])
    );

    PE u_pe11_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][8]),
        //Up part
        .weight_i(weight_i[185]),
        .sum_i(sum_o[10][9]),
        //Right part
        .data_o(data_o[11][9]),
        //Down part
        .sum_o(sum_o[11][9])
    );

    PE u_pe11_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][9]),
        //Up part
        .weight_i(weight_i[186]),
        .sum_i(sum_o[10][10]),
        //Right part
        .data_o(data_o[11][10]),
        //Down part
        .sum_o(sum_o[11][10])
    );

    PE u_pe11_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][10]),
        //Up part
        .weight_i(weight_i[187]),
        .sum_i(sum_o[10][11]),
        //Right part
        .data_o(data_o[11][11]),
        //Down part
        .sum_o(sum_o[11][11])
    );

    PE u_pe11_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][11]),
        //Up part
        .weight_i(weight_i[188]),
        .sum_i(sum_o[10][12]),
        //Right part
        .data_o(data_o[11][12]),
        //Down part
        .sum_o(sum_o[11][12])
    );

    PE u_pe11_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][12]),
        //Up part
        .weight_i(weight_i[189]),
        .sum_i(sum_o[10][13]),
        //Right part
        .data_o(data_o[11][13]),
        //Down part
        .sum_o(sum_o[11][13])
    );

    PE u_pe11_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][13]),
        //Up part
        .weight_i(weight_i[190]),
        .sum_i(sum_o[10][14]),
        //Right part
        .data_o(data_o[11][14]),
        //Down part
        .sum_o(sum_o[11][14])
    );

    PE u_pe11_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[11][14]),
        //Up part
        .weight_i(weight_i[191]),
        .sum_i(sum_o[10][15]),
        //Right part
        .data_o(data_o[11][15]),
        //Down part
        .sum_o(sum_o[11][15])
    );

    //'12'th row
    PE u_pe12_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[12]),
        //Up part
        .weight_i(weight_i[192]),
        .sum_i(sum_o[11][0]),
        //Right part
        .data_o(data_o[12][0]),
        //Down part
        .sum_o(sum_o[12][0])
    );

    PE u_pe12_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][0]),
        //Up part
        .weight_i(weight_i[193]),
        .sum_i(sum_o[11][1]),
        //Right part
        .data_o(data_o[12][1]),
        //Down part
        .sum_o(sum_o[12][1])
    );

    PE u_pe12_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][1]),
        //Up part
        .weight_i(weight_i[194]),
        .sum_i(sum_o[11][2]),
        //Right part
        .data_o(data_o[12][2]),
        //Down part
        .sum_o(sum_o[12][2])
    );

    PE u_pe12_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][2]),
        //Up part
        .weight_i(weight_i[195]),
        .sum_i(sum_o[11][3]),
        //Right part
        .data_o(data_o[12][3]),
        //Down part
        .sum_o(sum_o[12][3])
    );

    PE u_pe12_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][3]),
        //Up part
        .weight_i(weight_i[196]),
        .sum_i(sum_o[11][4]),
        //Right part
        .data_o(data_o[12][4]),
        //Down part
        .sum_o(sum_o[12][4])
    );

    PE u_pe12_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][4]),
        //Up part
        .weight_i(weight_i[197]),
        .sum_i(sum_o[11][5]),
        //Right part
        .data_o(data_o[12][5]),
        //Down part
        .sum_o(sum_o[12][5])
    );

    PE u_pe12_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][5]),
        //Up part
        .weight_i(weight_i[198]),
        .sum_i(sum_o[11][6]),
        //Right part
        .data_o(data_o[12][6]),
        //Down part
        .sum_o(sum_o[12][6])
    );

    PE u_pe12_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][6]),
        //Up part
        .weight_i(weight_i[199]),
        .sum_i(sum_o[11][7]),
        //Right part
        .data_o(data_o[12][7]),
        //Down part
        .sum_o(sum_o[12][7])
    );

    PE u_pe12_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][7]),
        //Up part
        .weight_i(weight_i[200]),
        .sum_i(sum_o[11][8]),
        //Right part
        .data_o(data_o[12][8]),
        //Down part
        .sum_o(sum_o[12][8])
    );

    PE u_pe12_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][8]),
        //Up part
        .weight_i(weight_i[201]),
        .sum_i(sum_o[11][9]),
        //Right part
        .data_o(data_o[12][9]),
        //Down part
        .sum_o(sum_o[12][9])
    );

    PE u_pe12_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][9]),
        //Up part
        .weight_i(weight_i[202]),
        .sum_i(sum_o[11][10]),
        //Right part
        .data_o(data_o[12][10]),
        //Down part
        .sum_o(sum_o[12][10])
    );

    PE u_pe12_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][10]),
        //Up part
        .weight_i(weight_i[203]),
        .sum_i(sum_o[11][11]),
        //Right part
        .data_o(data_o[12][11]),
        //Down part
        .sum_o(sum_o[12][11])
    );

    PE u_pe12_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][11]),
        //Up part
        .weight_i(weight_i[204]),
        .sum_i(sum_o[11][12]),
        //Right part
        .data_o(data_o[12][12]),
        //Down part
        .sum_o(sum_o[12][12])
    );

    PE u_pe12_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][12]),
        //Up part
        .weight_i(weight_i[205]),
        .sum_i(sum_o[11][13]),
        //Right part
        .data_o(data_o[12][13]),
        //Down part
        .sum_o(sum_o[12][13])
    );

    PE u_pe12_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][13]),
        //Up part
        .weight_i(weight_i[206]),
        .sum_i(sum_o[11][14]),
        //Right part
        .data_o(data_o[12][14]),
        //Down part
        .sum_o(sum_o[12][14])
    );

    PE u_pe12_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[12][14]),
        //Up part
        .weight_i(weight_i[207]),
        .sum_i(sum_o[11][15]),
        //Right part
        .data_o(data_o[12][15]),
        //Down part
        .sum_o(sum_o[12][15])
    );

    //'13'th row
    PE u_pe13_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[13]),
        //Up part
        .weight_i(weight_i[208]),
        .sum_i(sum_o[12][0]),
        //Right part
        .data_o(data_o[13][0]),
        //Down part
        .sum_o(sum_o[13][0])
    );

    PE u_pe13_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][0]),
        //Up part
        .weight_i(weight_i[209]),
        .sum_i(sum_o[12][1]),
        //Right part
        .data_o(data_o[13][1]),
        //Down part
        .sum_o(sum_o[13][1])
    );

    PE u_pe13_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][1]),
        //Up part
        .weight_i(weight_i[210]),
        .sum_i(sum_o[12][2]),
        //Right part
        .data_o(data_o[13][2]),
        //Down part
        .sum_o(sum_o[13][2])
    );

    PE u_pe13_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][2]),
        //Up part
        .weight_i(weight_i[211]),
        .sum_i(sum_o[12][3]),
        //Right part
        .data_o(data_o[13][3]),
        //Down part
        .sum_o(sum_o[13][3])
    );

    PE u_pe13_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][3]),
        //Up part
        .weight_i(weight_i[212]),
        .sum_i(sum_o[12][4]),
        //Right part
        .data_o(data_o[13][4]),
        //Down part
        .sum_o(sum_o[13][4])
    );

    PE u_pe13_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][4]),
        //Up part
        .weight_i(weight_i[213]),
        .sum_i(sum_o[12][5]),
        //Right part
        .data_o(data_o[13][5]),
        //Down part
        .sum_o(sum_o[13][5])
    );

    PE u_pe13_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][5]),
        //Up part
        .weight_i(weight_i[214]),
        .sum_i(sum_o[12][6]),
        //Right part
        .data_o(data_o[13][6]),
        //Down part
        .sum_o(sum_o[13][6])
    );

    PE u_pe13_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][6]),
        //Up part
        .weight_i(weight_i[215]),
        .sum_i(sum_o[12][7]),
        //Right part
        .data_o(data_o[13][7]),
        //Down part
        .sum_o(sum_o[13][7])
    );

    PE u_pe13_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][7]),
        //Up part
        .weight_i(weight_i[216]),
        .sum_i(sum_o[12][8]),
        //Right part
        .data_o(data_o[13][8]),
        //Down part
        .sum_o(sum_o[13][8])
    );

    PE u_pe13_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][8]),
        //Up part
        .weight_i(weight_i[217]),
        .sum_i(sum_o[12][9]),
        //Right part
        .data_o(data_o[13][9]),
        //Down part
        .sum_o(sum_o[13][9])
    );

    PE u_pe13_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][9]),
        //Up part
        .weight_i(weight_i[218]),
        .sum_i(sum_o[12][10]),
        //Right part
        .data_o(data_o[13][10]),
        //Down part
        .sum_o(sum_o[13][10])
    );

    PE u_pe13_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][10]),
        //Up part
        .weight_i(weight_i[219]),
        .sum_i(sum_o[12][11]),
        //Right part
        .data_o(data_o[13][11]),
        //Down part
        .sum_o(sum_o[13][11])
    );

    PE u_pe13_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][11]),
        //Up part
        .weight_i(weight_i[220]),
        .sum_i(sum_o[12][12]),
        //Right part
        .data_o(data_o[13][12]),
        //Down part
        .sum_o(sum_o[13][12])
    );

    PE u_pe13_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][12]),
        //Up part
        .weight_i(weight_i[221]),
        .sum_i(sum_o[12][13]),
        //Right part
        .data_o(data_o[13][13]),
        //Down part
        .sum_o(sum_o[13][13])
    );

    PE u_pe13_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][13]),
        //Up part
        .weight_i(weight_i[222]),
        .sum_i(sum_o[12][14]),
        //Right part
        .data_o(data_o[13][14]),
        //Down part
        .sum_o(sum_o[13][14])
    );

    PE u_pe13_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[13][14]),
        //Up part
        .weight_i(weight_i[223]),
        .sum_i(sum_o[12][15]),
        //Right part
        .data_o(data_o[13][15]),
        //Down part
        .sum_o(sum_o[13][15])
    );

    //'14'th row
    PE u_pe14_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[14]),
        //Up part
        .weight_i(weight_i[224]),
        .sum_i(sum_o[13][0]),
        //Right part
        .data_o(data_o[14][0]),
        //Down part
        .sum_o(sum_o[14][0])
    );

    PE u_pe14_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][0]),
        //Up part
        .weight_i(weight_i[225]),
        .sum_i(sum_o[13][1]),
        //Right part
        .data_o(data_o[14][1]),
        //Down part
        .sum_o(sum_o[14][1])
    );

    PE u_pe14_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][1]),
        //Up part
        .weight_i(weight_i[226]),
        .sum_i(sum_o[13][2]),
        //Right part
        .data_o(data_o[14][2]),
        //Down part
        .sum_o(sum_o[14][2])
    );

    PE u_pe14_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][2]),
        //Up part
        .weight_i(weight_i[227]),
        .sum_i(sum_o[13][3]),
        //Right part
        .data_o(data_o[14][3]),
        //Down part
        .sum_o(sum_o[14][3])
    );

    PE u_pe14_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][3]),
        //Up part
        .weight_i(weight_i[228]),
        .sum_i(sum_o[13][4]),
        //Right part
        .data_o(data_o[14][4]),
        //Down part
        .sum_o(sum_o[14][4])
    );

    PE u_pe14_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][4]),
        //Up part
        .weight_i(weight_i[229]),
        .sum_i(sum_o[13][5]),
        //Right part
        .data_o(data_o[14][5]),
        //Down part
        .sum_o(sum_o[14][5])
    );

    PE u_pe14_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][5]),
        //Up part
        .weight_i(weight_i[230]),
        .sum_i(sum_o[13][6]),
        //Right part
        .data_o(data_o[14][6]),
        //Down part
        .sum_o(sum_o[14][6])
    );

    PE u_pe14_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][6]),
        //Up part
        .weight_i(weight_i[231]),
        .sum_i(sum_o[13][7]),
        //Right part
        .data_o(data_o[14][7]),
        //Down part
        .sum_o(sum_o[14][7])
    );

    PE u_pe14_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][7]),
        //Up part
        .weight_i(weight_i[232]),
        .sum_i(sum_o[13][8]),
        //Right part
        .data_o(data_o[14][8]),
        //Down part
        .sum_o(sum_o[14][8])
    );

    PE u_pe14_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][8]),
        //Up part
        .weight_i(weight_i[233]),
        .sum_i(sum_o[13][9]),
        //Right part
        .data_o(data_o[14][9]),
        //Down part
        .sum_o(sum_o[14][9])
    );

    PE u_pe14_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][9]),
        //Up part
        .weight_i(weight_i[234]),
        .sum_i(sum_o[13][10]),
        //Right part
        .data_o(data_o[14][10]),
        //Down part
        .sum_o(sum_o[14][10])
    );

    PE u_pe14_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][10]),
        //Up part
        .weight_i(weight_i[235]),
        .sum_i(sum_o[13][11]),
        //Right part
        .data_o(data_o[14][11]),
        //Down part
        .sum_o(sum_o[14][11])
    );

    PE u_pe14_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][11]),
        //Up part
        .weight_i(weight_i[236]),
        .sum_i(sum_o[13][12]),
        //Right part
        .data_o(data_o[14][12]),
        //Down part
        .sum_o(sum_o[14][12])
    );

    PE u_pe14_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][12]),
        //Up part
        .weight_i(weight_i[237]),
        .sum_i(sum_o[13][13]),
        //Right part
        .data_o(data_o[14][13]),
        //Down part
        .sum_o(sum_o[14][13])
    );

    PE u_pe14_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][13]),
        //Up part
        .weight_i(weight_i[238]),
        .sum_i(sum_o[13][14]),
        //Right part
        .data_o(data_o[14][14]),
        //Down part
        .sum_o(sum_o[14][14])
    );

    PE u_pe14_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[14][14]),
        //Up part
        .weight_i(weight_i[239]),
        .sum_i(sum_o[13][15]),
        //Right part
        .data_o(data_o[14][15]),
        //Down part
        .sum_o(sum_o[14][15])
    );

    //'15'th row
    PE u_pe15_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[15]),
        //Up part
        .weight_i(weight_i[240]),
        .sum_i(sum_o[14][0]),
        //Right part
        .data_o(data_o[15][0]),
        //Down part
        .sum_o(sum_o[15][0])
    );

    PE u_pe15_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][0]),
        //Up part
        .weight_i(weight_i[241]),
        .sum_i(sum_o[14][1]),
        //Right part
        .data_o(data_o[15][1]),
        //Down part
        .sum_o(sum_o[15][1])
    );

    PE u_pe15_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][1]),
        //Up part
        .weight_i(weight_i[242]),
        .sum_i(sum_o[14][2]),
        //Right part
        .data_o(data_o[15][2]),
        //Down part
        .sum_o(sum_o[15][2])
    );

    PE u_pe15_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][2]),
        //Up part
        .weight_i(weight_i[243]),
        .sum_i(sum_o[14][3]),
        //Right part
        .data_o(data_o[15][3]),
        //Down part
        .sum_o(sum_o[15][3])
    );

    PE u_pe15_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][3]),
        //Up part
        .weight_i(weight_i[244]),
        .sum_i(sum_o[14][4]),
        //Right part
        .data_o(data_o[15][4]),
        //Down part
        .sum_o(sum_o[15][4])
    );

    PE u_pe15_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][4]),
        //Up part
        .weight_i(weight_i[245]),
        .sum_i(sum_o[14][5]),
        //Right part
        .data_o(data_o[15][5]),
        //Down part
        .sum_o(sum_o[15][5])
    );

    PE u_pe15_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][5]),
        //Up part
        .weight_i(weight_i[246]),
        .sum_i(sum_o[14][6]),
        //Right part
        .data_o(data_o[15][6]),
        //Down part
        .sum_o(sum_o[15][6])
    );

    PE u_pe15_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][6]),
        //Up part
        .weight_i(weight_i[247]),
        .sum_i(sum_o[14][7]),
        //Right part
        .data_o(data_o[15][7]),
        //Down part
        .sum_o(sum_o[15][7])
    );

    PE u_pe15_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][7]),
        //Up part
        .weight_i(weight_i[248]),
        .sum_i(sum_o[14][8]),
        //Right part
        .data_o(data_o[15][8]),
        //Down part
        .sum_o(sum_o[15][8])
    );

    PE u_pe15_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][8]),
        //Up part
        .weight_i(weight_i[249]),
        .sum_i(sum_o[14][9]),
        //Right part
        .data_o(data_o[15][9]),
        //Down part
        .sum_o(sum_o[15][9])
    );

    PE u_pe15_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][9]),
        //Up part
        .weight_i(weight_i[250]),
        .sum_i(sum_o[14][10]),
        //Right part
        .data_o(data_o[15][10]),
        //Down part
        .sum_o(sum_o[15][10])
    );

    PE u_pe15_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][10]),
        //Up part
        .weight_i(weight_i[251]),
        .sum_i(sum_o[14][11]),
        //Right part
        .data_o(data_o[15][11]),
        //Down part
        .sum_o(sum_o[15][11])
    );

    PE u_pe15_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][11]),
        //Up part
        .weight_i(weight_i[252]),
        .sum_i(sum_o[14][12]),
        //Right part
        .data_o(data_o[15][12]),
        //Down part
        .sum_o(sum_o[15][12])
    );

    PE u_pe15_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][12]),
        //Up part
        .weight_i(weight_i[253]),
        .sum_i(sum_o[14][13]),
        //Right part
        .data_o(data_o[15][13]),
        //Down part
        .sum_o(sum_o[15][13])
    );

    PE u_pe15_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][13]),
        //Up part
        .weight_i(weight_i[254]),
        .sum_i(sum_o[14][14]),
        //Right part
        .data_o(data_o[15][14]),
        //Down part
        .sum_o(sum_o[15][14])
    );

    PE u_pe15_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[15][14]),
        //Up part
        .weight_i(weight_i[255]),
        .sum_i(sum_o[14][15]),
        //Right part
        .data_o(data_o[15][15]),
        //Down part
        .sum_o(sum_o[15][15])
    );

    //'16'th row
    PE u_pe16_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[16]),
        //Up part
        .weight_i(weight_i[256]),
        .sum_i(sum_o[15][0]),
        //Right part
        .data_o(data_o[16][0]),
        //Down part
        .sum_o(sum_o[16][0])
    );

    PE u_pe16_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][0]),
        //Up part
        .weight_i(weight_i[257]),
        .sum_i(sum_o[15][1]),
        //Right part
        .data_o(data_o[16][1]),
        //Down part
        .sum_o(sum_o[16][1])
    );

    PE u_pe16_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][1]),
        //Up part
        .weight_i(weight_i[258]),
        .sum_i(sum_o[15][2]),
        //Right part
        .data_o(data_o[16][2]),
        //Down part
        .sum_o(sum_o[16][2])
    );

    PE u_pe16_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][2]),
        //Up part
        .weight_i(weight_i[259]),
        .sum_i(sum_o[15][3]),
        //Right part
        .data_o(data_o[16][3]),
        //Down part
        .sum_o(sum_o[16][3])
    );

    PE u_pe16_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][3]),
        //Up part
        .weight_i(weight_i[260]),
        .sum_i(sum_o[15][4]),
        //Right part
        .data_o(data_o[16][4]),
        //Down part
        .sum_o(sum_o[16][4])
    );

    PE u_pe16_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][4]),
        //Up part
        .weight_i(weight_i[261]),
        .sum_i(sum_o[15][5]),
        //Right part
        .data_o(data_o[16][5]),
        //Down part
        .sum_o(sum_o[16][5])
    );

    PE u_pe16_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][5]),
        //Up part
        .weight_i(weight_i[262]),
        .sum_i(sum_o[15][6]),
        //Right part
        .data_o(data_o[16][6]),
        //Down part
        .sum_o(sum_o[16][6])
    );

    PE u_pe16_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][6]),
        //Up part
        .weight_i(weight_i[263]),
        .sum_i(sum_o[15][7]),
        //Right part
        .data_o(data_o[16][7]),
        //Down part
        .sum_o(sum_o[16][7])
    );

    PE u_pe16_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][7]),
        //Up part
        .weight_i(weight_i[264]),
        .sum_i(sum_o[15][8]),
        //Right part
        .data_o(data_o[16][8]),
        //Down part
        .sum_o(sum_o[16][8])
    );

    PE u_pe16_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][8]),
        //Up part
        .weight_i(weight_i[265]),
        .sum_i(sum_o[15][9]),
        //Right part
        .data_o(data_o[16][9]),
        //Down part
        .sum_o(sum_o[16][9])
    );

    PE u_pe16_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][9]),
        //Up part
        .weight_i(weight_i[266]),
        .sum_i(sum_o[15][10]),
        //Right part
        .data_o(data_o[16][10]),
        //Down part
        .sum_o(sum_o[16][10])
    );

    PE u_pe16_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][10]),
        //Up part
        .weight_i(weight_i[267]),
        .sum_i(sum_o[15][11]),
        //Right part
        .data_o(data_o[16][11]),
        //Down part
        .sum_o(sum_o[16][11])
    );

    PE u_pe16_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][11]),
        //Up part
        .weight_i(weight_i[268]),
        .sum_i(sum_o[15][12]),
        //Right part
        .data_o(data_o[16][12]),
        //Down part
        .sum_o(sum_o[16][12])
    );

    PE u_pe16_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][12]),
        //Up part
        .weight_i(weight_i[269]),
        .sum_i(sum_o[15][13]),
        //Right part
        .data_o(data_o[16][13]),
        //Down part
        .sum_o(sum_o[16][13])
    );

    PE u_pe16_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][13]),
        //Up part
        .weight_i(weight_i[270]),
        .sum_i(sum_o[15][14]),
        //Right part
        .data_o(data_o[16][14]),
        //Down part
        .sum_o(sum_o[16][14])
    );

    PE u_pe16_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[16][14]),
        //Up part
        .weight_i(weight_i[271]),
        .sum_i(sum_o[15][15]),
        //Right part
        .data_o(data_o[16][15]),
        //Down part
        .sum_o(sum_o[16][15])
    );

    //'17'th row
    PE u_pe17_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[17]),
        //Up part
        .weight_i(weight_i[272]),
        .sum_i(sum_o[16][0]),
        //Right part
        .data_o(data_o[17][0]),
        //Down part
        .sum_o(sum_o[17][0])
    );

    PE u_pe17_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][0]),
        //Up part
        .weight_i(weight_i[273]),
        .sum_i(sum_o[16][1]),
        //Right part
        .data_o(data_o[17][1]),
        //Down part
        .sum_o(sum_o[17][1])
    );

    PE u_pe17_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][1]),
        //Up part
        .weight_i(weight_i[274]),
        .sum_i(sum_o[16][2]),
        //Right part
        .data_o(data_o[17][2]),
        //Down part
        .sum_o(sum_o[17][2])
    );

    PE u_pe17_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][2]),
        //Up part
        .weight_i(weight_i[275]),
        .sum_i(sum_o[16][3]),
        //Right part
        .data_o(data_o[17][3]),
        //Down part
        .sum_o(sum_o[17][3])
    );

    PE u_pe17_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][3]),
        //Up part
        .weight_i(weight_i[276]),
        .sum_i(sum_o[16][4]),
        //Right part
        .data_o(data_o[17][4]),
        //Down part
        .sum_o(sum_o[17][4])
    );

    PE u_pe17_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][4]),
        //Up part
        .weight_i(weight_i[277]),
        .sum_i(sum_o[16][5]),
        //Right part
        .data_o(data_o[17][5]),
        //Down part
        .sum_o(sum_o[17][5])
    );

    PE u_pe17_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][5]),
        //Up part
        .weight_i(weight_i[278]),
        .sum_i(sum_o[16][6]),
        //Right part
        .data_o(data_o[17][6]),
        //Down part
        .sum_o(sum_o[17][6])
    );

    PE u_pe17_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][6]),
        //Up part
        .weight_i(weight_i[279]),
        .sum_i(sum_o[16][7]),
        //Right part
        .data_o(data_o[17][7]),
        //Down part
        .sum_o(sum_o[17][7])
    );

    PE u_pe17_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][7]),
        //Up part
        .weight_i(weight_i[280]),
        .sum_i(sum_o[16][8]),
        //Right part
        .data_o(data_o[17][8]),
        //Down part
        .sum_o(sum_o[17][8])
    );

    PE u_pe17_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][8]),
        //Up part
        .weight_i(weight_i[281]),
        .sum_i(sum_o[16][9]),
        //Right part
        .data_o(data_o[17][9]),
        //Down part
        .sum_o(sum_o[17][9])
    );

    PE u_pe17_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][9]),
        //Up part
        .weight_i(weight_i[282]),
        .sum_i(sum_o[16][10]),
        //Right part
        .data_o(data_o[17][10]),
        //Down part
        .sum_o(sum_o[17][10])
    );

    PE u_pe17_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][10]),
        //Up part
        .weight_i(weight_i[283]),
        .sum_i(sum_o[16][11]),
        //Right part
        .data_o(data_o[17][11]),
        //Down part
        .sum_o(sum_o[17][11])
    );

    PE u_pe17_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][11]),
        //Up part
        .weight_i(weight_i[284]),
        .sum_i(sum_o[16][12]),
        //Right part
        .data_o(data_o[17][12]),
        //Down part
        .sum_o(sum_o[17][12])
    );

    PE u_pe17_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][12]),
        //Up part
        .weight_i(weight_i[285]),
        .sum_i(sum_o[16][13]),
        //Right part
        .data_o(data_o[17][13]),
        //Down part
        .sum_o(sum_o[17][13])
    );

    PE u_pe17_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][13]),
        //Up part
        .weight_i(weight_i[286]),
        .sum_i(sum_o[16][14]),
        //Right part
        .data_o(data_o[17][14]),
        //Down part
        .sum_o(sum_o[17][14])
    );

    PE u_pe17_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[17][14]),
        //Up part
        .weight_i(weight_i[287]),
        .sum_i(sum_o[16][15]),
        //Right part
        .data_o(data_o[17][15]),
        //Down part
        .sum_o(sum_o[17][15])
    );

    //'18'th row
    PE u_pe18_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[18]),
        //Up part
        .weight_i(weight_i[288]),
        .sum_i(sum_o[17][0]),
        //Right part
        .data_o(data_o[18][0]),
        //Down part
        .sum_o(sum_o[18][0])
    );

    PE u_pe18_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][0]),
        //Up part
        .weight_i(weight_i[289]),
        .sum_i(sum_o[17][1]),
        //Right part
        .data_o(data_o[18][1]),
        //Down part
        .sum_o(sum_o[18][1])
    );

    PE u_pe18_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][1]),
        //Up part
        .weight_i(weight_i[290]),
        .sum_i(sum_o[17][2]),
        //Right part
        .data_o(data_o[18][2]),
        //Down part
        .sum_o(sum_o[18][2])
    );

    PE u_pe18_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][2]),
        //Up part
        .weight_i(weight_i[291]),
        .sum_i(sum_o[17][3]),
        //Right part
        .data_o(data_o[18][3]),
        //Down part
        .sum_o(sum_o[18][3])
    );

    PE u_pe18_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][3]),
        //Up part
        .weight_i(weight_i[292]),
        .sum_i(sum_o[17][4]),
        //Right part
        .data_o(data_o[18][4]),
        //Down part
        .sum_o(sum_o[18][4])
    );

    PE u_pe18_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][4]),
        //Up part
        .weight_i(weight_i[293]),
        .sum_i(sum_o[17][5]),
        //Right part
        .data_o(data_o[18][5]),
        //Down part
        .sum_o(sum_o[18][5])
    );

    PE u_pe18_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][5]),
        //Up part
        .weight_i(weight_i[294]),
        .sum_i(sum_o[17][6]),
        //Right part
        .data_o(data_o[18][6]),
        //Down part
        .sum_o(sum_o[18][6])
    );

    PE u_pe18_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][6]),
        //Up part
        .weight_i(weight_i[295]),
        .sum_i(sum_o[17][7]),
        //Right part
        .data_o(data_o[18][7]),
        //Down part
        .sum_o(sum_o[18][7])
    );

    PE u_pe18_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][7]),
        //Up part
        .weight_i(weight_i[296]),
        .sum_i(sum_o[17][8]),
        //Right part
        .data_o(data_o[18][8]),
        //Down part
        .sum_o(sum_o[18][8])
    );

    PE u_pe18_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][8]),
        //Up part
        .weight_i(weight_i[297]),
        .sum_i(sum_o[17][9]),
        //Right part
        .data_o(data_o[18][9]),
        //Down part
        .sum_o(sum_o[18][9])
    );

    PE u_pe18_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][9]),
        //Up part
        .weight_i(weight_i[298]),
        .sum_i(sum_o[17][10]),
        //Right part
        .data_o(data_o[18][10]),
        //Down part
        .sum_o(sum_o[18][10])
    );

    PE u_pe18_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][10]),
        //Up part
        .weight_i(weight_i[299]),
        .sum_i(sum_o[17][11]),
        //Right part
        .data_o(data_o[18][11]),
        //Down part
        .sum_o(sum_o[18][11])
    );

    PE u_pe18_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][11]),
        //Up part
        .weight_i(weight_i[300]),
        .sum_i(sum_o[17][12]),
        //Right part
        .data_o(data_o[18][12]),
        //Down part
        .sum_o(sum_o[18][12])
    );

    PE u_pe18_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][12]),
        //Up part
        .weight_i(weight_i[301]),
        .sum_i(sum_o[17][13]),
        //Right part
        .data_o(data_o[18][13]),
        //Down part
        .sum_o(sum_o[18][13])
    );

    PE u_pe18_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][13]),
        //Up part
        .weight_i(weight_i[302]),
        .sum_i(sum_o[17][14]),
        //Right part
        .data_o(data_o[18][14]),
        //Down part
        .sum_o(sum_o[18][14])
    );

    PE u_pe18_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[18][14]),
        //Up part
        .weight_i(weight_i[303]),
        .sum_i(sum_o[17][15]),
        //Right part
        .data_o(data_o[18][15]),
        //Down part
        .sum_o(sum_o[18][15])
    );

    //'19'th row
    PE u_pe19_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[19]),
        //Up part
        .weight_i(weight_i[304]),
        .sum_i(sum_o[18][0]),
        //Right part
        .data_o(data_o[19][0]),
        //Down part
        .sum_o(sum_o[19][0])
    );

    PE u_pe19_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][0]),
        //Up part
        .weight_i(weight_i[305]),
        .sum_i(sum_o[18][1]),
        //Right part
        .data_o(data_o[19][1]),
        //Down part
        .sum_o(sum_o[19][1])
    );

    PE u_pe19_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][1]),
        //Up part
        .weight_i(weight_i[306]),
        .sum_i(sum_o[18][2]),
        //Right part
        .data_o(data_o[19][2]),
        //Down part
        .sum_o(sum_o[19][2])
    );

    PE u_pe19_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][2]),
        //Up part
        .weight_i(weight_i[307]),
        .sum_i(sum_o[18][3]),
        //Right part
        .data_o(data_o[19][3]),
        //Down part
        .sum_o(sum_o[19][3])
    );

    PE u_pe19_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][3]),
        //Up part
        .weight_i(weight_i[308]),
        .sum_i(sum_o[18][4]),
        //Right part
        .data_o(data_o[19][4]),
        //Down part
        .sum_o(sum_o[19][4])
    );

    PE u_pe19_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][4]),
        //Up part
        .weight_i(weight_i[309]),
        .sum_i(sum_o[18][5]),
        //Right part
        .data_o(data_o[19][5]),
        //Down part
        .sum_o(sum_o[19][5])
    );

    PE u_pe19_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][5]),
        //Up part
        .weight_i(weight_i[310]),
        .sum_i(sum_o[18][6]),
        //Right part
        .data_o(data_o[19][6]),
        //Down part
        .sum_o(sum_o[19][6])
    );

    PE u_pe19_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][6]),
        //Up part
        .weight_i(weight_i[311]),
        .sum_i(sum_o[18][7]),
        //Right part
        .data_o(data_o[19][7]),
        //Down part
        .sum_o(sum_o[19][7])
    );

    PE u_pe19_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][7]),
        //Up part
        .weight_i(weight_i[312]),
        .sum_i(sum_o[18][8]),
        //Right part
        .data_o(data_o[19][8]),
        //Down part
        .sum_o(sum_o[19][8])
    );

    PE u_pe19_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][8]),
        //Up part
        .weight_i(weight_i[313]),
        .sum_i(sum_o[18][9]),
        //Right part
        .data_o(data_o[19][9]),
        //Down part
        .sum_o(sum_o[19][9])
    );

    PE u_pe19_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][9]),
        //Up part
        .weight_i(weight_i[314]),
        .sum_i(sum_o[18][10]),
        //Right part
        .data_o(data_o[19][10]),
        //Down part
        .sum_o(sum_o[19][10])
    );

    PE u_pe19_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][10]),
        //Up part
        .weight_i(weight_i[315]),
        .sum_i(sum_o[18][11]),
        //Right part
        .data_o(data_o[19][11]),
        //Down part
        .sum_o(sum_o[19][11])
    );

    PE u_pe19_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][11]),
        //Up part
        .weight_i(weight_i[316]),
        .sum_i(sum_o[18][12]),
        //Right part
        .data_o(data_o[19][12]),
        //Down part
        .sum_o(sum_o[19][12])
    );

    PE u_pe19_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][12]),
        //Up part
        .weight_i(weight_i[317]),
        .sum_i(sum_o[18][13]),
        //Right part
        .data_o(data_o[19][13]),
        //Down part
        .sum_o(sum_o[19][13])
    );

    PE u_pe19_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][13]),
        //Up part
        .weight_i(weight_i[318]),
        .sum_i(sum_o[18][14]),
        //Right part
        .data_o(data_o[19][14]),
        //Down part
        .sum_o(sum_o[19][14])
    );

    PE u_pe19_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[19][14]),
        //Up part
        .weight_i(weight_i[319]),
        .sum_i(sum_o[18][15]),
        //Right part
        .data_o(data_o[19][15]),
        //Down part
        .sum_o(sum_o[19][15])
    );

    //'20'th row
    PE u_pe20_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[20]),
        //Up part
        .weight_i(weight_i[320]),
        .sum_i(sum_o[19][0]),
        //Right part
        .data_o(data_o[20][0]),
        //Down part
        .sum_o(sum_o[20][0])
    );

    PE u_pe20_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][0]),
        //Up part
        .weight_i(weight_i[321]),
        .sum_i(sum_o[19][1]),
        //Right part
        .data_o(data_o[20][1]),
        //Down part
        .sum_o(sum_o[20][1])
    );

    PE u_pe20_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][1]),
        //Up part
        .weight_i(weight_i[322]),
        .sum_i(sum_o[19][2]),
        //Right part
        .data_o(data_o[20][2]),
        //Down part
        .sum_o(sum_o[20][2])
    );

    PE u_pe20_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][2]),
        //Up part
        .weight_i(weight_i[323]),
        .sum_i(sum_o[19][3]),
        //Right part
        .data_o(data_o[20][3]),
        //Down part
        .sum_o(sum_o[20][3])
    );

    PE u_pe20_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][3]),
        //Up part
        .weight_i(weight_i[324]),
        .sum_i(sum_o[19][4]),
        //Right part
        .data_o(data_o[20][4]),
        //Down part
        .sum_o(sum_o[20][4])
    );

    PE u_pe20_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][4]),
        //Up part
        .weight_i(weight_i[325]),
        .sum_i(sum_o[19][5]),
        //Right part
        .data_o(data_o[20][5]),
        //Down part
        .sum_o(sum_o[20][5])
    );

    PE u_pe20_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][5]),
        //Up part
        .weight_i(weight_i[326]),
        .sum_i(sum_o[19][6]),
        //Right part
        .data_o(data_o[20][6]),
        //Down part
        .sum_o(sum_o[20][6])
    );

    PE u_pe20_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][6]),
        //Up part
        .weight_i(weight_i[327]),
        .sum_i(sum_o[19][7]),
        //Right part
        .data_o(data_o[20][7]),
        //Down part
        .sum_o(sum_o[20][7])
    );

    PE u_pe20_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][7]),
        //Up part
        .weight_i(weight_i[328]),
        .sum_i(sum_o[19][8]),
        //Right part
        .data_o(data_o[20][8]),
        //Down part
        .sum_o(sum_o[20][8])
    );

    PE u_pe20_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][8]),
        //Up part
        .weight_i(weight_i[329]),
        .sum_i(sum_o[19][9]),
        //Right part
        .data_o(data_o[20][9]),
        //Down part
        .sum_o(sum_o[20][9])
    );

    PE u_pe20_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][9]),
        //Up part
        .weight_i(weight_i[330]),
        .sum_i(sum_o[19][10]),
        //Right part
        .data_o(data_o[20][10]),
        //Down part
        .sum_o(sum_o[20][10])
    );

    PE u_pe20_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][10]),
        //Up part
        .weight_i(weight_i[331]),
        .sum_i(sum_o[19][11]),
        //Right part
        .data_o(data_o[20][11]),
        //Down part
        .sum_o(sum_o[20][11])
    );

    PE u_pe20_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][11]),
        //Up part
        .weight_i(weight_i[332]),
        .sum_i(sum_o[19][12]),
        //Right part
        .data_o(data_o[20][12]),
        //Down part
        .sum_o(sum_o[20][12])
    );

    PE u_pe20_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][12]),
        //Up part
        .weight_i(weight_i[333]),
        .sum_i(sum_o[19][13]),
        //Right part
        .data_o(data_o[20][13]),
        //Down part
        .sum_o(sum_o[20][13])
    );

    PE u_pe20_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][13]),
        //Up part
        .weight_i(weight_i[334]),
        .sum_i(sum_o[19][14]),
        //Right part
        .data_o(data_o[20][14]),
        //Down part
        .sum_o(sum_o[20][14])
    );

    PE u_pe20_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[20][14]),
        //Up part
        .weight_i(weight_i[335]),
        .sum_i(sum_o[19][15]),
        //Right part
        .data_o(data_o[20][15]),
        //Down part
        .sum_o(sum_o[20][15])
    );

    //'21'th row
    PE u_pe21_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[21]),
        //Up part
        .weight_i(weight_i[336]),
        .sum_i(sum_o[20][0]),
        //Right part
        .data_o(data_o[21][0]),
        //Down part
        .sum_o(sum_o[21][0])
    );

    PE u_pe21_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][0]),
        //Up part
        .weight_i(weight_i[337]),
        .sum_i(sum_o[20][1]),
        //Right part
        .data_o(data_o[21][1]),
        //Down part
        .sum_o(sum_o[21][1])
    );

    PE u_pe21_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][1]),
        //Up part
        .weight_i(weight_i[338]),
        .sum_i(sum_o[20][2]),
        //Right part
        .data_o(data_o[21][2]),
        //Down part
        .sum_o(sum_o[21][2])
    );

    PE u_pe21_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][2]),
        //Up part
        .weight_i(weight_i[339]),
        .sum_i(sum_o[20][3]),
        //Right part
        .data_o(data_o[21][3]),
        //Down part
        .sum_o(sum_o[21][3])
    );

    PE u_pe21_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][3]),
        //Up part
        .weight_i(weight_i[340]),
        .sum_i(sum_o[20][4]),
        //Right part
        .data_o(data_o[21][4]),
        //Down part
        .sum_o(sum_o[21][4])
    );

    PE u_pe21_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][4]),
        //Up part
        .weight_i(weight_i[341]),
        .sum_i(sum_o[20][5]),
        //Right part
        .data_o(data_o[21][5]),
        //Down part
        .sum_o(sum_o[21][5])
    );

    PE u_pe21_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][5]),
        //Up part
        .weight_i(weight_i[342]),
        .sum_i(sum_o[20][6]),
        //Right part
        .data_o(data_o[21][6]),
        //Down part
        .sum_o(sum_o[21][6])
    );

    PE u_pe21_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][6]),
        //Up part
        .weight_i(weight_i[343]),
        .sum_i(sum_o[20][7]),
        //Right part
        .data_o(data_o[21][7]),
        //Down part
        .sum_o(sum_o[21][7])
    );

    PE u_pe21_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][7]),
        //Up part
        .weight_i(weight_i[344]),
        .sum_i(sum_o[20][8]),
        //Right part
        .data_o(data_o[21][8]),
        //Down part
        .sum_o(sum_o[21][8])
    );

    PE u_pe21_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][8]),
        //Up part
        .weight_i(weight_i[345]),
        .sum_i(sum_o[20][9]),
        //Right part
        .data_o(data_o[21][9]),
        //Down part
        .sum_o(sum_o[21][9])
    );

    PE u_pe21_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][9]),
        //Up part
        .weight_i(weight_i[346]),
        .sum_i(sum_o[20][10]),
        //Right part
        .data_o(data_o[21][10]),
        //Down part
        .sum_o(sum_o[21][10])
    );

    PE u_pe21_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][10]),
        //Up part
        .weight_i(weight_i[347]),
        .sum_i(sum_o[20][11]),
        //Right part
        .data_o(data_o[21][11]),
        //Down part
        .sum_o(sum_o[21][11])
    );

    PE u_pe21_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][11]),
        //Up part
        .weight_i(weight_i[348]),
        .sum_i(sum_o[20][12]),
        //Right part
        .data_o(data_o[21][12]),
        //Down part
        .sum_o(sum_o[21][12])
    );

    PE u_pe21_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][12]),
        //Up part
        .weight_i(weight_i[349]),
        .sum_i(sum_o[20][13]),
        //Right part
        .data_o(data_o[21][13]),
        //Down part
        .sum_o(sum_o[21][13])
    );

    PE u_pe21_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][13]),
        //Up part
        .weight_i(weight_i[350]),
        .sum_i(sum_o[20][14]),
        //Right part
        .data_o(data_o[21][14]),
        //Down part
        .sum_o(sum_o[21][14])
    );

    PE u_pe21_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[21][14]),
        //Up part
        .weight_i(weight_i[351]),
        .sum_i(sum_o[20][15]),
        //Right part
        .data_o(data_o[21][15]),
        //Down part
        .sum_o(sum_o[21][15])
    );

    //'22'th row
    PE u_pe22_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[22]),
        //Up part
        .weight_i(weight_i[352]),
        .sum_i(sum_o[21][0]),
        //Right part
        .data_o(data_o[22][0]),
        //Down part
        .sum_o(sum_o[22][0])
    );

    PE u_pe22_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][0]),
        //Up part
        .weight_i(weight_i[353]),
        .sum_i(sum_o[21][1]),
        //Right part
        .data_o(data_o[22][1]),
        //Down part
        .sum_o(sum_o[22][1])
    );

    PE u_pe22_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][1]),
        //Up part
        .weight_i(weight_i[354]),
        .sum_i(sum_o[21][2]),
        //Right part
        .data_o(data_o[22][2]),
        //Down part
        .sum_o(sum_o[22][2])
    );

    PE u_pe22_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][2]),
        //Up part
        .weight_i(weight_i[355]),
        .sum_i(sum_o[21][3]),
        //Right part
        .data_o(data_o[22][3]),
        //Down part
        .sum_o(sum_o[22][3])
    );

    PE u_pe22_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][3]),
        //Up part
        .weight_i(weight_i[356]),
        .sum_i(sum_o[21][4]),
        //Right part
        .data_o(data_o[22][4]),
        //Down part
        .sum_o(sum_o[22][4])
    );

    PE u_pe22_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][4]),
        //Up part
        .weight_i(weight_i[357]),
        .sum_i(sum_o[21][5]),
        //Right part
        .data_o(data_o[22][5]),
        //Down part
        .sum_o(sum_o[22][5])
    );

    PE u_pe22_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][5]),
        //Up part
        .weight_i(weight_i[358]),
        .sum_i(sum_o[21][6]),
        //Right part
        .data_o(data_o[22][6]),
        //Down part
        .sum_o(sum_o[22][6])
    );

    PE u_pe22_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][6]),
        //Up part
        .weight_i(weight_i[359]),
        .sum_i(sum_o[21][7]),
        //Right part
        .data_o(data_o[22][7]),
        //Down part
        .sum_o(sum_o[22][7])
    );

    PE u_pe22_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][7]),
        //Up part
        .weight_i(weight_i[360]),
        .sum_i(sum_o[21][8]),
        //Right part
        .data_o(data_o[22][8]),
        //Down part
        .sum_o(sum_o[22][8])
    );

    PE u_pe22_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][8]),
        //Up part
        .weight_i(weight_i[361]),
        .sum_i(sum_o[21][9]),
        //Right part
        .data_o(data_o[22][9]),
        //Down part
        .sum_o(sum_o[22][9])
    );

    PE u_pe22_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][9]),
        //Up part
        .weight_i(weight_i[362]),
        .sum_i(sum_o[21][10]),
        //Right part
        .data_o(data_o[22][10]),
        //Down part
        .sum_o(sum_o[22][10])
    );

    PE u_pe22_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][10]),
        //Up part
        .weight_i(weight_i[363]),
        .sum_i(sum_o[21][11]),
        //Right part
        .data_o(data_o[22][11]),
        //Down part
        .sum_o(sum_o[22][11])
    );

    PE u_pe22_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][11]),
        //Up part
        .weight_i(weight_i[364]),
        .sum_i(sum_o[21][12]),
        //Right part
        .data_o(data_o[22][12]),
        //Down part
        .sum_o(sum_o[22][12])
    );

    PE u_pe22_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][12]),
        //Up part
        .weight_i(weight_i[365]),
        .sum_i(sum_o[21][13]),
        //Right part
        .data_o(data_o[22][13]),
        //Down part
        .sum_o(sum_o[22][13])
    );

    PE u_pe22_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][13]),
        //Up part
        .weight_i(weight_i[366]),
        .sum_i(sum_o[21][14]),
        //Right part
        .data_o(data_o[22][14]),
        //Down part
        .sum_o(sum_o[22][14])
    );

    PE u_pe22_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[22][14]),
        //Up part
        .weight_i(weight_i[367]),
        .sum_i(sum_o[21][15]),
        //Right part
        .data_o(data_o[22][15]),
        //Down part
        .sum_o(sum_o[22][15])
    );

    //'23'th row
    PE u_pe23_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[23]),
        //Up part
        .weight_i(weight_i[368]),
        .sum_i(sum_o[22][0]),
        //Right part
        .data_o(data_o[23][0]),
        //Down part
        .sum_o(sum_o[23][0])
    );

    PE u_pe23_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][0]),
        //Up part
        .weight_i(weight_i[369]),
        .sum_i(sum_o[22][1]),
        //Right part
        .data_o(data_o[23][1]),
        //Down part
        .sum_o(sum_o[23][1])
    );

    PE u_pe23_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][1]),
        //Up part
        .weight_i(weight_i[370]),
        .sum_i(sum_o[22][2]),
        //Right part
        .data_o(data_o[23][2]),
        //Down part
        .sum_o(sum_o[23][2])
    );

    PE u_pe23_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][2]),
        //Up part
        .weight_i(weight_i[371]),
        .sum_i(sum_o[22][3]),
        //Right part
        .data_o(data_o[23][3]),
        //Down part
        .sum_o(sum_o[23][3])
    );

    PE u_pe23_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][3]),
        //Up part
        .weight_i(weight_i[372]),
        .sum_i(sum_o[22][4]),
        //Right part
        .data_o(data_o[23][4]),
        //Down part
        .sum_o(sum_o[23][4])
    );

    PE u_pe23_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][4]),
        //Up part
        .weight_i(weight_i[373]),
        .sum_i(sum_o[22][5]),
        //Right part
        .data_o(data_o[23][5]),
        //Down part
        .sum_o(sum_o[23][5])
    );

    PE u_pe23_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][5]),
        //Up part
        .weight_i(weight_i[374]),
        .sum_i(sum_o[22][6]),
        //Right part
        .data_o(data_o[23][6]),
        //Down part
        .sum_o(sum_o[23][6])
    );

    PE u_pe23_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][6]),
        //Up part
        .weight_i(weight_i[375]),
        .sum_i(sum_o[22][7]),
        //Right part
        .data_o(data_o[23][7]),
        //Down part
        .sum_o(sum_o[23][7])
    );

    PE u_pe23_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][7]),
        //Up part
        .weight_i(weight_i[376]),
        .sum_i(sum_o[22][8]),
        //Right part
        .data_o(data_o[23][8]),
        //Down part
        .sum_o(sum_o[23][8])
    );

    PE u_pe23_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][8]),
        //Up part
        .weight_i(weight_i[377]),
        .sum_i(sum_o[22][9]),
        //Right part
        .data_o(data_o[23][9]),
        //Down part
        .sum_o(sum_o[23][9])
    );

    PE u_pe23_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][9]),
        //Up part
        .weight_i(weight_i[378]),
        .sum_i(sum_o[22][10]),
        //Right part
        .data_o(data_o[23][10]),
        //Down part
        .sum_o(sum_o[23][10])
    );

    PE u_pe23_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][10]),
        //Up part
        .weight_i(weight_i[379]),
        .sum_i(sum_o[22][11]),
        //Right part
        .data_o(data_o[23][11]),
        //Down part
        .sum_o(sum_o[23][11])
    );

    PE u_pe23_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][11]),
        //Up part
        .weight_i(weight_i[380]),
        .sum_i(sum_o[22][12]),
        //Right part
        .data_o(data_o[23][12]),
        //Down part
        .sum_o(sum_o[23][12])
    );

    PE u_pe23_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][12]),
        //Up part
        .weight_i(weight_i[381]),
        .sum_i(sum_o[22][13]),
        //Right part
        .data_o(data_o[23][13]),
        //Down part
        .sum_o(sum_o[23][13])
    );

    PE u_pe23_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][13]),
        //Up part
        .weight_i(weight_i[382]),
        .sum_i(sum_o[22][14]),
        //Right part
        .data_o(data_o[23][14]),
        //Down part
        .sum_o(sum_o[23][14])
    );

    PE u_pe23_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[23][14]),
        //Up part
        .weight_i(weight_i[383]),
        .sum_i(sum_o[22][15]),
        //Right part
        .data_o(data_o[23][15]),
        //Down part
        .sum_o(sum_o[23][15])
    );

    //'24'th row
    PE u_pe24_0(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_i[24]),
        //Up part
        .weight_i(weight_i[384]),
        .sum_i(sum_o[23][0]),
        //Right part
        .data_o(data_o[24][0]),
        //Down part
        .sum_o(sum_o[24][0])
    );

    PE u_pe24_1(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][0]),
        //Up part
        .weight_i(weight_i[385]),
        .sum_i(sum_o[23][1]),
        //Right part
        .data_o(data_o[24][1]),
        //Down part
        .sum_o(sum_o[24][1])
    );

    PE u_pe24_2(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][1]),
        //Up part
        .weight_i(weight_i[386]),
        .sum_i(sum_o[23][2]),
        //Right part
        .data_o(data_o[24][2]),
        //Down part
        .sum_o(sum_o[24][2])
    );

    PE u_pe24_3(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][2]),
        //Up part
        .weight_i(weight_i[387]),
        .sum_i(sum_o[23][3]),
        //Right part
        .data_o(data_o[24][3]),
        //Down part
        .sum_o(sum_o[24][3])
    );

    PE u_pe24_4(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][3]),
        //Up part
        .weight_i(weight_i[388]),
        .sum_i(sum_o[23][4]),
        //Right part
        .data_o(data_o[24][4]),
        //Down part
        .sum_o(sum_o[24][4])
    );

    PE u_pe24_5(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][4]),
        //Up part
        .weight_i(weight_i[389]),
        .sum_i(sum_o[23][5]),
        //Right part
        .data_o(data_o[24][5]),
        //Down part
        .sum_o(sum_o[24][5])
    );

    PE u_pe24_6(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][5]),
        //Up part
        .weight_i(weight_i[390]),
        .sum_i(sum_o[23][6]),
        //Right part
        .data_o(data_o[24][6]),
        //Down part
        .sum_o(sum_o[24][6])
    );

    PE u_pe24_7(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][6]),
        //Up part
        .weight_i(weight_i[391]),
        .sum_i(sum_o[23][7]),
        //Right part
        .data_o(data_o[24][7]),
        //Down part
        .sum_o(sum_o[24][7])
    );

    PE u_pe24_8(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][7]),
        //Up part
        .weight_i(weight_i[392]),
        .sum_i(sum_o[23][8]),
        //Right part
        .data_o(data_o[24][8]),
        //Down part
        .sum_o(sum_o[24][8])
    );

    PE u_pe24_9(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][8]),
        //Up part
        .weight_i(weight_i[393]),
        .sum_i(sum_o[23][9]),
        //Right part
        .data_o(data_o[24][9]),
        //Down part
        .sum_o(sum_o[24][9])
    );

    PE u_pe24_10(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][9]),
        //Up part
        .weight_i(weight_i[394]),
        .sum_i(sum_o[23][10]),
        //Right part
        .data_o(data_o[24][10]),
        //Down part
        .sum_o(sum_o[24][10])
    );

    PE u_pe24_11(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][10]),
        //Up part
        .weight_i(weight_i[395]),
        .sum_i(sum_o[23][11]),
        //Right part
        .data_o(data_o[24][11]),
        //Down part
        .sum_o(sum_o[24][11])
    );

    PE u_pe24_12(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][11]),
        //Up part
        .weight_i(weight_i[396]),
        .sum_i(sum_o[23][12]),
        //Right part
        .data_o(data_o[24][12]),
        //Down part
        .sum_o(sum_o[24][12])
    );

    PE u_pe24_13(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][12]),
        //Up part
        .weight_i(weight_i[397]),
        .sum_i(sum_o[23][13]),
        //Right part
        .data_o(data_o[24][13]),
        //Down part
        .sum_o(sum_o[24][13])
    );

    PE u_pe24_14(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][13]),
        //Up part
        .weight_i(weight_i[398]),
        .sum_i(sum_o[23][14]),
        //Right part
        .data_o(data_o[24][14]),
        //Down part
        .sum_o(sum_o[24][14])
    );

    PE u_pe24_15(
        .clk(clk),
        .rst_n(rst_n),
        //Left part
        .data_i(data_o[24][14]),
        //Up part
        .weight_i(weight_i[399]),
        .sum_i(sum_o[23][15]),
        //Right part
        .data_o(data_o[24][15]),
        //Down part
        .sum_o(sum_o[24][15])
    );



    always_ff @(posedge clk) begin


    end

    always_comb begin

    end


endmodule