//version 2022-01-19
//editor IM SUHYEOK

module SA_ctrl
(
    input   wire                        clk,
    input   wire                        rst_n,
    input   wire                        start_i,        
    input   wire                        data_last_i,
    input   wire                        [1:0] nth_conv_i,
    input   wire                        conv_done_i,
    output  wire                        data_enable_o,          //data setup
    output  wire                        weight_start_o,         //weight buffer
    output  wire                        weight_stop_o           //SA
);

    localparam          S_IDLE      = 2'd0,
                        S_CONV      = 2'd1,
                        S_CONV_N    = 2'd2,
                        S_CONV2_N   = 2'd3;

    reg                 [1:0] state, state_n;
    reg                 data_enable;
    reg                 [4:0] cnt, cnt_n;
    reg                 weight_start;
    reg                 weight_stop;


    always_ff @(posedge clk) begin
        if(!rst_n) begin
            state <= S_IDLE;
            cnt <= 5'd0;
        end
        else begin
            state <= state_n;
            cnt <= cnt_n;
        end
    end

    always_comb begin
        data_enable = 1'b0;
        weight_start = 1'b0;
        state_n = state;
        cnt_n   = cnt;

        case(state)
            S_IDLE: begin
                weight_stop = 1'b0;
                if(start_i) begin
                    state_n = S_CONV;
                    weight_start = 1'b1;
                end
            end
            S_CONV: begin
                cnt_n = cnt + 'd1;
                if(cnt < 'd27) begin
                    weight_stop = 1'b0;
                end
                else begin
                    weight_stop = 1'b1;
                end

                if(cnt == 'd26) begin
                    weight_start = 1'b0;
                end

                if(cnt == 'd28) begin
                    cnt_n = 'd0;
                    data_enable = 1'b1;
                    if (nth_conv_i == 0) begin
                        state_n = S_CONV_N;
                    end 
                    else begin
                        state_n = S_CONV2_N;
                    end
                end
            end
            S_CONV_N: begin
                data_enable = 1'b1;
                if(conv_done_i) begin
                    data_enable = 1'b0;
                    state_n = S_IDLE;
                end
            end
            S_CONV2_N : begin
                if(!conv_done_i) begin
                    data_enable = 1'b1;
                    if(data_last_i) begin
                        data_enable = 1'b0;
                        state_n = S_CONV;
                    end
                end
                else begin
                    data_enable = 1'b0;
                    state_n = S_IDLE;
                end
            end    
        endcase
    end

    assign data_enable_o        = data_enable;
    assign weight_stop_o        = weight_stop;
    assign weight_start_o       = weight_start;

endmodule